// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 11 2025 23:51:26

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_g,
    T01,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_g;
    output T01;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__50432;
    wire N__50431;
    wire N__50430;
    wire N__50421;
    wire N__50420;
    wire N__50419;
    wire N__50412;
    wire N__50411;
    wire N__50410;
    wire N__50403;
    wire N__50402;
    wire N__50401;
    wire N__50394;
    wire N__50393;
    wire N__50392;
    wire N__50385;
    wire N__50384;
    wire N__50383;
    wire N__50376;
    wire N__50375;
    wire N__50374;
    wire N__50367;
    wire N__50366;
    wire N__50365;
    wire N__50358;
    wire N__50357;
    wire N__50356;
    wire N__50349;
    wire N__50348;
    wire N__50347;
    wire N__50340;
    wire N__50339;
    wire N__50338;
    wire N__50331;
    wire N__50330;
    wire N__50329;
    wire N__50322;
    wire N__50321;
    wire N__50320;
    wire N__50313;
    wire N__50312;
    wire N__50311;
    wire N__50304;
    wire N__50303;
    wire N__50302;
    wire N__50295;
    wire N__50294;
    wire N__50293;
    wire N__50286;
    wire N__50285;
    wire N__50284;
    wire N__50267;
    wire N__50264;
    wire N__50261;
    wire N__50260;
    wire N__50259;
    wire N__50258;
    wire N__50255;
    wire N__50252;
    wire N__50249;
    wire N__50246;
    wire N__50237;
    wire N__50236;
    wire N__50235;
    wire N__50232;
    wire N__50229;
    wire N__50226;
    wire N__50223;
    wire N__50220;
    wire N__50213;
    wire N__50212;
    wire N__50209;
    wire N__50206;
    wire N__50201;
    wire N__50198;
    wire N__50197;
    wire N__50194;
    wire N__50193;
    wire N__50190;
    wire N__50187;
    wire N__50184;
    wire N__50177;
    wire N__50174;
    wire N__50173;
    wire N__50172;
    wire N__50169;
    wire N__50166;
    wire N__50163;
    wire N__50162;
    wire N__50157;
    wire N__50154;
    wire N__50151;
    wire N__50144;
    wire N__50143;
    wire N__50138;
    wire N__50135;
    wire N__50134;
    wire N__50133;
    wire N__50132;
    wire N__50129;
    wire N__50126;
    wire N__50121;
    wire N__50118;
    wire N__50115;
    wire N__50108;
    wire N__50105;
    wire N__50102;
    wire N__50101;
    wire N__50100;
    wire N__50099;
    wire N__50098;
    wire N__50095;
    wire N__50092;
    wire N__50089;
    wire N__50084;
    wire N__50079;
    wire N__50074;
    wire N__50071;
    wire N__50066;
    wire N__50063;
    wire N__50062;
    wire N__50059;
    wire N__50056;
    wire N__50055;
    wire N__50054;
    wire N__50053;
    wire N__50052;
    wire N__50051;
    wire N__50050;
    wire N__50049;
    wire N__50048;
    wire N__50047;
    wire N__50042;
    wire N__50035;
    wire N__50034;
    wire N__50033;
    wire N__50032;
    wire N__50031;
    wire N__50028;
    wire N__50027;
    wire N__50018;
    wire N__50015;
    wire N__50010;
    wire N__50007;
    wire N__50006;
    wire N__50005;
    wire N__50002;
    wire N__50001;
    wire N__50000;
    wire N__49999;
    wire N__49998;
    wire N__49995;
    wire N__49994;
    wire N__49991;
    wire N__49990;
    wire N__49987;
    wire N__49984;
    wire N__49983;
    wire N__49982;
    wire N__49981;
    wire N__49980;
    wire N__49979;
    wire N__49978;
    wire N__49977;
    wire N__49976;
    wire N__49975;
    wire N__49970;
    wire N__49965;
    wire N__49964;
    wire N__49963;
    wire N__49962;
    wire N__49961;
    wire N__49960;
    wire N__49959;
    wire N__49958;
    wire N__49957;
    wire N__49956;
    wire N__49955;
    wire N__49954;
    wire N__49953;
    wire N__49952;
    wire N__49949;
    wire N__49946;
    wire N__49943;
    wire N__49934;
    wire N__49931;
    wire N__49928;
    wire N__49925;
    wire N__49922;
    wire N__49917;
    wire N__49914;
    wire N__49911;
    wire N__49902;
    wire N__49895;
    wire N__49890;
    wire N__49881;
    wire N__49872;
    wire N__49863;
    wire N__49860;
    wire N__49855;
    wire N__49852;
    wire N__49849;
    wire N__49846;
    wire N__49837;
    wire N__49834;
    wire N__49831;
    wire N__49818;
    wire N__49815;
    wire N__49810;
    wire N__49801;
    wire N__49798;
    wire N__49795;
    wire N__49790;
    wire N__49787;
    wire N__49778;
    wire N__49777;
    wire N__49774;
    wire N__49773;
    wire N__49770;
    wire N__49769;
    wire N__49766;
    wire N__49763;
    wire N__49760;
    wire N__49757;
    wire N__49754;
    wire N__49749;
    wire N__49742;
    wire N__49741;
    wire N__49738;
    wire N__49735;
    wire N__49734;
    wire N__49731;
    wire N__49728;
    wire N__49725;
    wire N__49720;
    wire N__49715;
    wire N__49714;
    wire N__49713;
    wire N__49710;
    wire N__49709;
    wire N__49706;
    wire N__49703;
    wire N__49700;
    wire N__49697;
    wire N__49694;
    wire N__49691;
    wire N__49688;
    wire N__49685;
    wire N__49682;
    wire N__49679;
    wire N__49674;
    wire N__49667;
    wire N__49666;
    wire N__49663;
    wire N__49660;
    wire N__49659;
    wire N__49656;
    wire N__49653;
    wire N__49650;
    wire N__49645;
    wire N__49640;
    wire N__49639;
    wire N__49638;
    wire N__49637;
    wire N__49636;
    wire N__49635;
    wire N__49632;
    wire N__49631;
    wire N__49630;
    wire N__49629;
    wire N__49628;
    wire N__49627;
    wire N__49626;
    wire N__49625;
    wire N__49624;
    wire N__49623;
    wire N__49620;
    wire N__49619;
    wire N__49618;
    wire N__49617;
    wire N__49616;
    wire N__49615;
    wire N__49614;
    wire N__49613;
    wire N__49604;
    wire N__49601;
    wire N__49594;
    wire N__49593;
    wire N__49592;
    wire N__49591;
    wire N__49590;
    wire N__49589;
    wire N__49588;
    wire N__49587;
    wire N__49586;
    wire N__49585;
    wire N__49584;
    wire N__49583;
    wire N__49582;
    wire N__49581;
    wire N__49580;
    wire N__49579;
    wire N__49578;
    wire N__49577;
    wire N__49576;
    wire N__49575;
    wire N__49574;
    wire N__49573;
    wire N__49572;
    wire N__49571;
    wire N__49570;
    wire N__49569;
    wire N__49568;
    wire N__49567;
    wire N__49556;
    wire N__49555;
    wire N__49554;
    wire N__49551;
    wire N__49550;
    wire N__49549;
    wire N__49548;
    wire N__49547;
    wire N__49546;
    wire N__49543;
    wire N__49538;
    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49532;
    wire N__49531;
    wire N__49530;
    wire N__49527;
    wire N__49520;
    wire N__49517;
    wire N__49512;
    wire N__49509;
    wire N__49498;
    wire N__49489;
    wire N__49482;
    wire N__49481;
    wire N__49480;
    wire N__49479;
    wire N__49476;
    wire N__49473;
    wire N__49470;
    wire N__49469;
    wire N__49466;
    wire N__49459;
    wire N__49458;
    wire N__49457;
    wire N__49456;
    wire N__49455;
    wire N__49454;
    wire N__49453;
    wire N__49452;
    wire N__49447;
    wire N__49436;
    wire N__49433;
    wire N__49430;
    wire N__49429;
    wire N__49426;
    wire N__49425;
    wire N__49424;
    wire N__49423;
    wire N__49422;
    wire N__49421;
    wire N__49420;
    wire N__49419;
    wire N__49418;
    wire N__49415;
    wire N__49408;
    wire N__49403;
    wire N__49400;
    wire N__49395;
    wire N__49392;
    wire N__49383;
    wire N__49372;
    wire N__49367;
    wire N__49364;
    wire N__49357;
    wire N__49354;
    wire N__49353;
    wire N__49352;
    wire N__49351;
    wire N__49350;
    wire N__49343;
    wire N__49340;
    wire N__49337;
    wire N__49336;
    wire N__49335;
    wire N__49334;
    wire N__49329;
    wire N__49322;
    wire N__49321;
    wire N__49320;
    wire N__49319;
    wire N__49318;
    wire N__49313;
    wire N__49304;
    wire N__49301;
    wire N__49298;
    wire N__49295;
    wire N__49288;
    wire N__49281;
    wire N__49278;
    wire N__49267;
    wire N__49264;
    wire N__49257;
    wire N__49250;
    wire N__49247;
    wire N__49242;
    wire N__49239;
    wire N__49232;
    wire N__49229;
    wire N__49224;
    wire N__49219;
    wire N__49210;
    wire N__49203;
    wire N__49196;
    wire N__49189;
    wire N__49182;
    wire N__49157;
    wire N__49154;
    wire N__49151;
    wire N__49148;
    wire N__49147;
    wire N__49146;
    wire N__49145;
    wire N__49144;
    wire N__49143;
    wire N__49142;
    wire N__49141;
    wire N__49140;
    wire N__49139;
    wire N__49138;
    wire N__49137;
    wire N__49136;
    wire N__49135;
    wire N__49134;
    wire N__49133;
    wire N__49132;
    wire N__49131;
    wire N__49130;
    wire N__49129;
    wire N__49128;
    wire N__49127;
    wire N__49126;
    wire N__49125;
    wire N__49124;
    wire N__49123;
    wire N__49122;
    wire N__49121;
    wire N__49120;
    wire N__49119;
    wire N__49118;
    wire N__49117;
    wire N__49116;
    wire N__49115;
    wire N__49114;
    wire N__49113;
    wire N__49112;
    wire N__49111;
    wire N__49110;
    wire N__49109;
    wire N__49108;
    wire N__49107;
    wire N__49106;
    wire N__49105;
    wire N__49104;
    wire N__49103;
    wire N__49102;
    wire N__49101;
    wire N__49100;
    wire N__49099;
    wire N__49098;
    wire N__49097;
    wire N__49096;
    wire N__49095;
    wire N__49094;
    wire N__49093;
    wire N__49092;
    wire N__49091;
    wire N__49090;
    wire N__49089;
    wire N__49088;
    wire N__49087;
    wire N__49086;
    wire N__49085;
    wire N__49084;
    wire N__49083;
    wire N__49082;
    wire N__49081;
    wire N__49080;
    wire N__49079;
    wire N__49078;
    wire N__49077;
    wire N__49076;
    wire N__49075;
    wire N__49074;
    wire N__49073;
    wire N__49072;
    wire N__49071;
    wire N__49070;
    wire N__49069;
    wire N__49068;
    wire N__49067;
    wire N__49066;
    wire N__49065;
    wire N__49064;
    wire N__49063;
    wire N__49062;
    wire N__49061;
    wire N__49060;
    wire N__49059;
    wire N__49058;
    wire N__49057;
    wire N__49056;
    wire N__49055;
    wire N__49054;
    wire N__49053;
    wire N__49052;
    wire N__49051;
    wire N__49050;
    wire N__49049;
    wire N__49048;
    wire N__49047;
    wire N__49046;
    wire N__49045;
    wire N__49044;
    wire N__49043;
    wire N__49042;
    wire N__49041;
    wire N__49040;
    wire N__49039;
    wire N__49038;
    wire N__49037;
    wire N__49036;
    wire N__49035;
    wire N__49034;
    wire N__49033;
    wire N__49032;
    wire N__49031;
    wire N__49030;
    wire N__49029;
    wire N__49028;
    wire N__49027;
    wire N__49026;
    wire N__49025;
    wire N__49024;
    wire N__49023;
    wire N__49022;
    wire N__49021;
    wire N__49020;
    wire N__49019;
    wire N__49018;
    wire N__49017;
    wire N__49016;
    wire N__49015;
    wire N__49014;
    wire N__49013;
    wire N__49012;
    wire N__49011;
    wire N__49010;
    wire N__49009;
    wire N__49008;
    wire N__48725;
    wire N__48722;
    wire N__48721;
    wire N__48720;
    wire N__48719;
    wire N__48718;
    wire N__48717;
    wire N__48716;
    wire N__48715;
    wire N__48714;
    wire N__48713;
    wire N__48712;
    wire N__48689;
    wire N__48686;
    wire N__48683;
    wire N__48682;
    wire N__48681;
    wire N__48680;
    wire N__48677;
    wire N__48674;
    wire N__48671;
    wire N__48668;
    wire N__48665;
    wire N__48662;
    wire N__48659;
    wire N__48658;
    wire N__48657;
    wire N__48656;
    wire N__48655;
    wire N__48654;
    wire N__48653;
    wire N__48652;
    wire N__48651;
    wire N__48650;
    wire N__48649;
    wire N__48648;
    wire N__48647;
    wire N__48646;
    wire N__48645;
    wire N__48644;
    wire N__48643;
    wire N__48642;
    wire N__48641;
    wire N__48640;
    wire N__48639;
    wire N__48638;
    wire N__48637;
    wire N__48636;
    wire N__48635;
    wire N__48634;
    wire N__48633;
    wire N__48632;
    wire N__48631;
    wire N__48630;
    wire N__48629;
    wire N__48628;
    wire N__48627;
    wire N__48626;
    wire N__48625;
    wire N__48624;
    wire N__48623;
    wire N__48622;
    wire N__48621;
    wire N__48620;
    wire N__48619;
    wire N__48618;
    wire N__48617;
    wire N__48616;
    wire N__48615;
    wire N__48614;
    wire N__48613;
    wire N__48612;
    wire N__48611;
    wire N__48610;
    wire N__48609;
    wire N__48608;
    wire N__48607;
    wire N__48606;
    wire N__48605;
    wire N__48604;
    wire N__48603;
    wire N__48602;
    wire N__48601;
    wire N__48600;
    wire N__48599;
    wire N__48598;
    wire N__48597;
    wire N__48596;
    wire N__48595;
    wire N__48594;
    wire N__48593;
    wire N__48592;
    wire N__48591;
    wire N__48590;
    wire N__48589;
    wire N__48588;
    wire N__48587;
    wire N__48586;
    wire N__48585;
    wire N__48584;
    wire N__48583;
    wire N__48582;
    wire N__48581;
    wire N__48580;
    wire N__48579;
    wire N__48578;
    wire N__48577;
    wire N__48576;
    wire N__48575;
    wire N__48574;
    wire N__48573;
    wire N__48572;
    wire N__48571;
    wire N__48570;
    wire N__48569;
    wire N__48568;
    wire N__48567;
    wire N__48566;
    wire N__48565;
    wire N__48564;
    wire N__48563;
    wire N__48560;
    wire N__48559;
    wire N__48558;
    wire N__48557;
    wire N__48556;
    wire N__48555;
    wire N__48554;
    wire N__48553;
    wire N__48552;
    wire N__48551;
    wire N__48550;
    wire N__48549;
    wire N__48548;
    wire N__48547;
    wire N__48546;
    wire N__48545;
    wire N__48544;
    wire N__48543;
    wire N__48542;
    wire N__48541;
    wire N__48540;
    wire N__48539;
    wire N__48538;
    wire N__48537;
    wire N__48536;
    wire N__48535;
    wire N__48534;
    wire N__48533;
    wire N__48532;
    wire N__48531;
    wire N__48530;
    wire N__48529;
    wire N__48528;
    wire N__48527;
    wire N__48526;
    wire N__48525;
    wire N__48524;
    wire N__48523;
    wire N__48522;
    wire N__48521;
    wire N__48520;
    wire N__48519;
    wire N__48518;
    wire N__48517;
    wire N__48516;
    wire N__48227;
    wire N__48224;
    wire N__48221;
    wire N__48218;
    wire N__48215;
    wire N__48214;
    wire N__48211;
    wire N__48208;
    wire N__48203;
    wire N__48200;
    wire N__48199;
    wire N__48194;
    wire N__48191;
    wire N__48188;
    wire N__48185;
    wire N__48182;
    wire N__48179;
    wire N__48178;
    wire N__48173;
    wire N__48172;
    wire N__48169;
    wire N__48168;
    wire N__48165;
    wire N__48162;
    wire N__48159;
    wire N__48152;
    wire N__48149;
    wire N__48148;
    wire N__48147;
    wire N__48144;
    wire N__48143;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48126;
    wire N__48121;
    wire N__48118;
    wire N__48113;
    wire N__48112;
    wire N__48111;
    wire N__48108;
    wire N__48107;
    wire N__48104;
    wire N__48101;
    wire N__48098;
    wire N__48095;
    wire N__48092;
    wire N__48087;
    wire N__48084;
    wire N__48079;
    wire N__48074;
    wire N__48073;
    wire N__48072;
    wire N__48067;
    wire N__48066;
    wire N__48063;
    wire N__48060;
    wire N__48057;
    wire N__48054;
    wire N__48049;
    wire N__48044;
    wire N__48041;
    wire N__48038;
    wire N__48035;
    wire N__48032;
    wire N__48029;
    wire N__48026;
    wire N__48023;
    wire N__48020;
    wire N__48017;
    wire N__48014;
    wire N__48011;
    wire N__48008;
    wire N__48005;
    wire N__48004;
    wire N__48003;
    wire N__48000;
    wire N__47995;
    wire N__47990;
    wire N__47989;
    wire N__47988;
    wire N__47985;
    wire N__47980;
    wire N__47975;
    wire N__47972;
    wire N__47969;
    wire N__47966;
    wire N__47963;
    wire N__47960;
    wire N__47959;
    wire N__47958;
    wire N__47955;
    wire N__47952;
    wire N__47949;
    wire N__47948;
    wire N__47945;
    wire N__47942;
    wire N__47939;
    wire N__47936;
    wire N__47931;
    wire N__47928;
    wire N__47925;
    wire N__47918;
    wire N__47915;
    wire N__47914;
    wire N__47913;
    wire N__47910;
    wire N__47907;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47891;
    wire N__47890;
    wire N__47887;
    wire N__47886;
    wire N__47885;
    wire N__47882;
    wire N__47879;
    wire N__47876;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47864;
    wire N__47861;
    wire N__47852;
    wire N__47851;
    wire N__47850;
    wire N__47845;
    wire N__47844;
    wire N__47841;
    wire N__47838;
    wire N__47835;
    wire N__47832;
    wire N__47829;
    wire N__47826;
    wire N__47823;
    wire N__47820;
    wire N__47817;
    wire N__47810;
    wire N__47809;
    wire N__47808;
    wire N__47805;
    wire N__47802;
    wire N__47801;
    wire N__47798;
    wire N__47793;
    wire N__47790;
    wire N__47787;
    wire N__47784;
    wire N__47781;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47765;
    wire N__47764;
    wire N__47761;
    wire N__47758;
    wire N__47757;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47745;
    wire N__47738;
    wire N__47735;
    wire N__47732;
    wire N__47729;
    wire N__47726;
    wire N__47723;
    wire N__47722;
    wire N__47717;
    wire N__47714;
    wire N__47711;
    wire N__47708;
    wire N__47707;
    wire N__47704;
    wire N__47703;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47687;
    wire N__47686;
    wire N__47683;
    wire N__47680;
    wire N__47679;
    wire N__47678;
    wire N__47675;
    wire N__47672;
    wire N__47669;
    wire N__47666;
    wire N__47663;
    wire N__47658;
    wire N__47655;
    wire N__47648;
    wire N__47647;
    wire N__47642;
    wire N__47639;
    wire N__47636;
    wire N__47635;
    wire N__47632;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47622;
    wire N__47615;
    wire N__47612;
    wire N__47609;
    wire N__47606;
    wire N__47603;
    wire N__47600;
    wire N__47599;
    wire N__47596;
    wire N__47595;
    wire N__47592;
    wire N__47589;
    wire N__47586;
    wire N__47579;
    wire N__47578;
    wire N__47573;
    wire N__47570;
    wire N__47569;
    wire N__47564;
    wire N__47561;
    wire N__47558;
    wire N__47555;
    wire N__47552;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47542;
    wire N__47541;
    wire N__47538;
    wire N__47533;
    wire N__47528;
    wire N__47527;
    wire N__47524;
    wire N__47523;
    wire N__47520;
    wire N__47515;
    wire N__47510;
    wire N__47507;
    wire N__47504;
    wire N__47501;
    wire N__47500;
    wire N__47497;
    wire N__47494;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47479;
    wire N__47474;
    wire N__47471;
    wire N__47470;
    wire N__47465;
    wire N__47462;
    wire N__47459;
    wire N__47456;
    wire N__47453;
    wire N__47452;
    wire N__47449;
    wire N__47446;
    wire N__47445;
    wire N__47440;
    wire N__47437;
    wire N__47434;
    wire N__47429;
    wire N__47426;
    wire N__47425;
    wire N__47422;
    wire N__47419;
    wire N__47418;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47402;
    wire N__47399;
    wire N__47396;
    wire N__47393;
    wire N__47392;
    wire N__47389;
    wire N__47386;
    wire N__47381;
    wire N__47378;
    wire N__47377;
    wire N__47376;
    wire N__47373;
    wire N__47368;
    wire N__47365;
    wire N__47362;
    wire N__47357;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47345;
    wire N__47344;
    wire N__47339;
    wire N__47336;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47324;
    wire N__47321;
    wire N__47318;
    wire N__47315;
    wire N__47312;
    wire N__47311;
    wire N__47310;
    wire N__47305;
    wire N__47302;
    wire N__47299;
    wire N__47294;
    wire N__47293;
    wire N__47290;
    wire N__47287;
    wire N__47286;
    wire N__47281;
    wire N__47278;
    wire N__47275;
    wire N__47270;
    wire N__47267;
    wire N__47264;
    wire N__47261;
    wire N__47258;
    wire N__47255;
    wire N__47254;
    wire N__47251;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47234;
    wire N__47231;
    wire N__47228;
    wire N__47227;
    wire N__47226;
    wire N__47225;
    wire N__47222;
    wire N__47219;
    wire N__47214;
    wire N__47207;
    wire N__47204;
    wire N__47201;
    wire N__47198;
    wire N__47195;
    wire N__47192;
    wire N__47191;
    wire N__47190;
    wire N__47187;
    wire N__47184;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47168;
    wire N__47167;
    wire N__47166;
    wire N__47165;
    wire N__47164;
    wire N__47163;
    wire N__47162;
    wire N__47161;
    wire N__47144;
    wire N__47141;
    wire N__47138;
    wire N__47135;
    wire N__47134;
    wire N__47131;
    wire N__47128;
    wire N__47125;
    wire N__47122;
    wire N__47121;
    wire N__47118;
    wire N__47115;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47103;
    wire N__47096;
    wire N__47095;
    wire N__47094;
    wire N__47091;
    wire N__47090;
    wire N__47087;
    wire N__47084;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47066;
    wire N__47063;
    wire N__47060;
    wire N__47053;
    wire N__47048;
    wire N__47045;
    wire N__47042;
    wire N__47041;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47028;
    wire N__47025;
    wire N__47018;
    wire N__47015;
    wire N__47012;
    wire N__47009;
    wire N__47006;
    wire N__47003;
    wire N__47000;
    wire N__46997;
    wire N__46996;
    wire N__46993;
    wire N__46990;
    wire N__46985;
    wire N__46982;
    wire N__46981;
    wire N__46976;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46966;
    wire N__46961;
    wire N__46960;
    wire N__46957;
    wire N__46954;
    wire N__46949;
    wire N__46948;
    wire N__46945;
    wire N__46942;
    wire N__46939;
    wire N__46934;
    wire N__46933;
    wire N__46928;
    wire N__46925;
    wire N__46922;
    wire N__46919;
    wire N__46916;
    wire N__46913;
    wire N__46910;
    wire N__46907;
    wire N__46906;
    wire N__46903;
    wire N__46900;
    wire N__46895;
    wire N__46892;
    wire N__46889;
    wire N__46886;
    wire N__46885;
    wire N__46880;
    wire N__46879;
    wire N__46876;
    wire N__46873;
    wire N__46870;
    wire N__46865;
    wire N__46862;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46854;
    wire N__46851;
    wire N__46848;
    wire N__46845;
    wire N__46840;
    wire N__46837;
    wire N__46836;
    wire N__46833;
    wire N__46830;
    wire N__46827;
    wire N__46820;
    wire N__46817;
    wire N__46816;
    wire N__46811;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46801;
    wire N__46796;
    wire N__46795;
    wire N__46792;
    wire N__46789;
    wire N__46786;
    wire N__46783;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46772;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46754;
    wire N__46751;
    wire N__46750;
    wire N__46747;
    wire N__46744;
    wire N__46739;
    wire N__46738;
    wire N__46735;
    wire N__46732;
    wire N__46729;
    wire N__46724;
    wire N__46721;
    wire N__46720;
    wire N__46717;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46698;
    wire N__46697;
    wire N__46694;
    wire N__46691;
    wire N__46688;
    wire N__46685;
    wire N__46676;
    wire N__46673;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46661;
    wire N__46660;
    wire N__46657;
    wire N__46654;
    wire N__46651;
    wire N__46646;
    wire N__46645;
    wire N__46642;
    wire N__46641;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46629;
    wire N__46624;
    wire N__46623;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46607;
    wire N__46604;
    wire N__46601;
    wire N__46598;
    wire N__46597;
    wire N__46594;
    wire N__46591;
    wire N__46590;
    wire N__46585;
    wire N__46582;
    wire N__46579;
    wire N__46574;
    wire N__46571;
    wire N__46570;
    wire N__46567;
    wire N__46564;
    wire N__46563;
    wire N__46562;
    wire N__46559;
    wire N__46554;
    wire N__46551;
    wire N__46544;
    wire N__46541;
    wire N__46538;
    wire N__46535;
    wire N__46532;
    wire N__46529;
    wire N__46528;
    wire N__46525;
    wire N__46522;
    wire N__46521;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46505;
    wire N__46502;
    wire N__46501;
    wire N__46498;
    wire N__46497;
    wire N__46494;
    wire N__46491;
    wire N__46488;
    wire N__46485;
    wire N__46482;
    wire N__46479;
    wire N__46478;
    wire N__46475;
    wire N__46472;
    wire N__46469;
    wire N__46466;
    wire N__46457;
    wire N__46454;
    wire N__46451;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46436;
    wire N__46433;
    wire N__46432;
    wire N__46431;
    wire N__46428;
    wire N__46425;
    wire N__46422;
    wire N__46417;
    wire N__46412;
    wire N__46409;
    wire N__46408;
    wire N__46407;
    wire N__46406;
    wire N__46403;
    wire N__46398;
    wire N__46395;
    wire N__46392;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46376;
    wire N__46373;
    wire N__46370;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46355;
    wire N__46352;
    wire N__46351;
    wire N__46348;
    wire N__46345;
    wire N__46344;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46328;
    wire N__46325;
    wire N__46324;
    wire N__46321;
    wire N__46320;
    wire N__46317;
    wire N__46314;
    wire N__46311;
    wire N__46308;
    wire N__46303;
    wire N__46302;
    wire N__46299;
    wire N__46296;
    wire N__46293;
    wire N__46286;
    wire N__46283;
    wire N__46280;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46272;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46256;
    wire N__46253;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46245;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46229;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46217;
    wire N__46214;
    wire N__46213;
    wire N__46208;
    wire N__46207;
    wire N__46204;
    wire N__46201;
    wire N__46198;
    wire N__46193;
    wire N__46190;
    wire N__46187;
    wire N__46184;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46162;
    wire N__46159;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46142;
    wire N__46139;
    wire N__46136;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46128;
    wire N__46123;
    wire N__46120;
    wire N__46117;
    wire N__46112;
    wire N__46111;
    wire N__46108;
    wire N__46105;
    wire N__46102;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46094;
    wire N__46091;
    wire N__46088;
    wire N__46085;
    wire N__46082;
    wire N__46079;
    wire N__46072;
    wire N__46067;
    wire N__46064;
    wire N__46063;
    wire N__46060;
    wire N__46057;
    wire N__46052;
    wire N__46051;
    wire N__46048;
    wire N__46045;
    wire N__46042;
    wire N__46037;
    wire N__46036;
    wire N__46035;
    wire N__46032;
    wire N__46029;
    wire N__46028;
    wire N__46025;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46009;
    wire N__46004;
    wire N__46001;
    wire N__45998;
    wire N__45995;
    wire N__45994;
    wire N__45991;
    wire N__45988;
    wire N__45987;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45971;
    wire N__45968;
    wire N__45967;
    wire N__45964;
    wire N__45963;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45951;
    wire N__45946;
    wire N__45945;
    wire N__45942;
    wire N__45939;
    wire N__45936;
    wire N__45929;
    wire N__45926;
    wire N__45923;
    wire N__45920;
    wire N__45919;
    wire N__45916;
    wire N__45913;
    wire N__45912;
    wire N__45907;
    wire N__45904;
    wire N__45901;
    wire N__45896;
    wire N__45895;
    wire N__45892;
    wire N__45891;
    wire N__45888;
    wire N__45885;
    wire N__45882;
    wire N__45877;
    wire N__45874;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45857;
    wire N__45854;
    wire N__45851;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45843;
    wire N__45838;
    wire N__45835;
    wire N__45832;
    wire N__45827;
    wire N__45824;
    wire N__45823;
    wire N__45820;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45800;
    wire N__45797;
    wire N__45794;
    wire N__45791;
    wire N__45788;
    wire N__45779;
    wire N__45776;
    wire N__45773;
    wire N__45772;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45762;
    wire N__45757;
    wire N__45752;
    wire N__45749;
    wire N__45748;
    wire N__45747;
    wire N__45740;
    wire N__45739;
    wire N__45736;
    wire N__45733;
    wire N__45728;
    wire N__45725;
    wire N__45722;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45714;
    wire N__45709;
    wire N__45706;
    wire N__45703;
    wire N__45698;
    wire N__45695;
    wire N__45694;
    wire N__45691;
    wire N__45688;
    wire N__45687;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45655;
    wire N__45650;
    wire N__45647;
    wire N__45646;
    wire N__45641;
    wire N__45640;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45626;
    wire N__45623;
    wire N__45622;
    wire N__45621;
    wire N__45620;
    wire N__45617;
    wire N__45612;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45592;
    wire N__45587;
    wire N__45584;
    wire N__45583;
    wire N__45578;
    wire N__45577;
    wire N__45574;
    wire N__45571;
    wire N__45568;
    wire N__45563;
    wire N__45562;
    wire N__45559;
    wire N__45556;
    wire N__45553;
    wire N__45550;
    wire N__45549;
    wire N__45548;
    wire N__45545;
    wire N__45542;
    wire N__45539;
    wire N__45536;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45509;
    wire N__45506;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45494;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45484;
    wire N__45479;
    wire N__45478;
    wire N__45477;
    wire N__45476;
    wire N__45471;
    wire N__45468;
    wire N__45465;
    wire N__45462;
    wire N__45459;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45443;
    wire N__45440;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45426;
    wire N__45423;
    wire N__45420;
    wire N__45417;
    wire N__45414;
    wire N__45411;
    wire N__45404;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45384;
    wire N__45379;
    wire N__45376;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45359;
    wire N__45356;
    wire N__45353;
    wire N__45352;
    wire N__45349;
    wire N__45346;
    wire N__45345;
    wire N__45342;
    wire N__45339;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45323;
    wire N__45322;
    wire N__45319;
    wire N__45316;
    wire N__45313;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45303;
    wire N__45298;
    wire N__45295;
    wire N__45294;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45278;
    wire N__45275;
    wire N__45272;
    wire N__45271;
    wire N__45268;
    wire N__45265;
    wire N__45264;
    wire N__45259;
    wire N__45256;
    wire N__45253;
    wire N__45248;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45232;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45222;
    wire N__45221;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45209;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45186;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45170;
    wire N__45169;
    wire N__45166;
    wire N__45163;
    wire N__45160;
    wire N__45157;
    wire N__45152;
    wire N__45151;
    wire N__45148;
    wire N__45145;
    wire N__45144;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45132;
    wire N__45127;
    wire N__45122;
    wire N__45119;
    wire N__45116;
    wire N__45113;
    wire N__45110;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45098;
    wire N__45097;
    wire N__45096;
    wire N__45095;
    wire N__45094;
    wire N__45093;
    wire N__45092;
    wire N__45091;
    wire N__45090;
    wire N__45089;
    wire N__45088;
    wire N__45087;
    wire N__45084;
    wire N__45083;
    wire N__45080;
    wire N__45079;
    wire N__45076;
    wire N__45075;
    wire N__45072;
    wire N__45071;
    wire N__45068;
    wire N__45067;
    wire N__45064;
    wire N__45063;
    wire N__45060;
    wire N__45059;
    wire N__45058;
    wire N__45055;
    wire N__45054;
    wire N__45051;
    wire N__45050;
    wire N__45047;
    wire N__45046;
    wire N__45045;
    wire N__45044;
    wire N__45041;
    wire N__45040;
    wire N__45039;
    wire N__45038;
    wire N__45037;
    wire N__45036;
    wire N__45021;
    wire N__45004;
    wire N__44989;
    wire N__44988;
    wire N__44987;
    wire N__44986;
    wire N__44985;
    wire N__44984;
    wire N__44983;
    wire N__44982;
    wire N__44981;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44969;
    wire N__44966;
    wire N__44965;
    wire N__44962;
    wire N__44961;
    wire N__44958;
    wire N__44957;
    wire N__44954;
    wire N__44953;
    wire N__44950;
    wire N__44945;
    wire N__44942;
    wire N__44935;
    wire N__44926;
    wire N__44925;
    wire N__44924;
    wire N__44921;
    wire N__44914;
    wire N__44897;
    wire N__44892;
    wire N__44891;
    wire N__44890;
    wire N__44883;
    wire N__44880;
    wire N__44879;
    wire N__44878;
    wire N__44877;
    wire N__44876;
    wire N__44875;
    wire N__44874;
    wire N__44873;
    wire N__44872;
    wire N__44869;
    wire N__44868;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44838;
    wire N__44829;
    wire N__44822;
    wire N__44819;
    wire N__44816;
    wire N__44809;
    wire N__44800;
    wire N__44797;
    wire N__44794;
    wire N__44789;
    wire N__44786;
    wire N__44783;
    wire N__44774;
    wire N__44771;
    wire N__44768;
    wire N__44765;
    wire N__44762;
    wire N__44759;
    wire N__44758;
    wire N__44757;
    wire N__44756;
    wire N__44755;
    wire N__44754;
    wire N__44753;
    wire N__44752;
    wire N__44747;
    wire N__44736;
    wire N__44735;
    wire N__44734;
    wire N__44733;
    wire N__44732;
    wire N__44731;
    wire N__44730;
    wire N__44729;
    wire N__44728;
    wire N__44727;
    wire N__44726;
    wire N__44725;
    wire N__44724;
    wire N__44723;
    wire N__44722;
    wire N__44721;
    wire N__44720;
    wire N__44719;
    wire N__44718;
    wire N__44717;
    wire N__44716;
    wire N__44715;
    wire N__44714;
    wire N__44713;
    wire N__44712;
    wire N__44711;
    wire N__44710;
    wire N__44709;
    wire N__44708;
    wire N__44707;
    wire N__44706;
    wire N__44705;
    wire N__44704;
    wire N__44701;
    wire N__44696;
    wire N__44679;
    wire N__44678;
    wire N__44677;
    wire N__44674;
    wire N__44669;
    wire N__44668;
    wire N__44667;
    wire N__44666;
    wire N__44665;
    wire N__44664;
    wire N__44663;
    wire N__44662;
    wire N__44661;
    wire N__44660;
    wire N__44659;
    wire N__44658;
    wire N__44657;
    wire N__44642;
    wire N__44625;
    wire N__44624;
    wire N__44623;
    wire N__44622;
    wire N__44621;
    wire N__44620;
    wire N__44609;
    wire N__44606;
    wire N__44599;
    wire N__44598;
    wire N__44597;
    wire N__44596;
    wire N__44595;
    wire N__44594;
    wire N__44593;
    wire N__44592;
    wire N__44591;
    wire N__44586;
    wire N__44581;
    wire N__44564;
    wire N__44557;
    wire N__44556;
    wire N__44553;
    wire N__44552;
    wire N__44551;
    wire N__44550;
    wire N__44545;
    wire N__44534;
    wire N__44527;
    wire N__44510;
    wire N__44507;
    wire N__44500;
    wire N__44489;
    wire N__44474;
    wire N__44471;
    wire N__44470;
    wire N__44469;
    wire N__44468;
    wire N__44467;
    wire N__44466;
    wire N__44465;
    wire N__44464;
    wire N__44463;
    wire N__44462;
    wire N__44461;
    wire N__44456;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44430;
    wire N__44429;
    wire N__44428;
    wire N__44427;
    wire N__44426;
    wire N__44421;
    wire N__44418;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44393;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44371;
    wire N__44366;
    wire N__44363;
    wire N__44362;
    wire N__44357;
    wire N__44356;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44339;
    wire N__44336;
    wire N__44335;
    wire N__44332;
    wire N__44329;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44309;
    wire N__44306;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44288;
    wire N__44285;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44269;
    wire N__44264;
    wire N__44261;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44249;
    wire N__44248;
    wire N__44245;
    wire N__44242;
    wire N__44239;
    wire N__44234;
    wire N__44231;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44223;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44205;
    wire N__44202;
    wire N__44199;
    wire N__44196;
    wire N__44191;
    wire N__44186;
    wire N__44183;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44171;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44156;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44138;
    wire N__44137;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44124;
    wire N__44119;
    wire N__44114;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44099;
    wire N__44096;
    wire N__44093;
    wire N__44090;
    wire N__44087;
    wire N__44084;
    wire N__44081;
    wire N__44078;
    wire N__44075;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44057;
    wire N__44054;
    wire N__44051;
    wire N__44048;
    wire N__44045;
    wire N__44042;
    wire N__44039;
    wire N__44036;
    wire N__44033;
    wire N__44030;
    wire N__44027;
    wire N__44024;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44012;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43985;
    wire N__43982;
    wire N__43979;
    wire N__43976;
    wire N__43973;
    wire N__43970;
    wire N__43967;
    wire N__43964;
    wire N__43961;
    wire N__43958;
    wire N__43955;
    wire N__43952;
    wire N__43949;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43937;
    wire N__43934;
    wire N__43931;
    wire N__43928;
    wire N__43925;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43901;
    wire N__43898;
    wire N__43895;
    wire N__43894;
    wire N__43893;
    wire N__43892;
    wire N__43889;
    wire N__43884;
    wire N__43881;
    wire N__43874;
    wire N__43873;
    wire N__43870;
    wire N__43867;
    wire N__43866;
    wire N__43863;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43841;
    wire N__43840;
    wire N__43837;
    wire N__43836;
    wire N__43833;
    wire N__43830;
    wire N__43827;
    wire N__43820;
    wire N__43817;
    wire N__43814;
    wire N__43811;
    wire N__43808;
    wire N__43807;
    wire N__43804;
    wire N__43801;
    wire N__43800;
    wire N__43799;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43789;
    wire N__43784;
    wire N__43781;
    wire N__43772;
    wire N__43769;
    wire N__43766;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43751;
    wire N__43748;
    wire N__43745;
    wire N__43742;
    wire N__43739;
    wire N__43736;
    wire N__43735;
    wire N__43734;
    wire N__43731;
    wire N__43728;
    wire N__43727;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43709;
    wire N__43706;
    wire N__43703;
    wire N__43700;
    wire N__43699;
    wire N__43698;
    wire N__43691;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43676;
    wire N__43673;
    wire N__43670;
    wire N__43667;
    wire N__43664;
    wire N__43661;
    wire N__43660;
    wire N__43659;
    wire N__43656;
    wire N__43651;
    wire N__43646;
    wire N__43643;
    wire N__43642;
    wire N__43641;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43594;
    wire N__43589;
    wire N__43586;
    wire N__43585;
    wire N__43584;
    wire N__43583;
    wire N__43580;
    wire N__43577;
    wire N__43574;
    wire N__43571;
    wire N__43562;
    wire N__43559;
    wire N__43558;
    wire N__43555;
    wire N__43554;
    wire N__43551;
    wire N__43548;
    wire N__43545;
    wire N__43538;
    wire N__43537;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43525;
    wire N__43524;
    wire N__43521;
    wire N__43516;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43499;
    wire N__43498;
    wire N__43497;
    wire N__43494;
    wire N__43489;
    wire N__43486;
    wire N__43483;
    wire N__43482;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43466;
    wire N__43463;
    wire N__43462;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43450;
    wire N__43445;
    wire N__43442;
    wire N__43441;
    wire N__43440;
    wire N__43437;
    wire N__43434;
    wire N__43429;
    wire N__43424;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43393;
    wire N__43388;
    wire N__43385;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43370;
    wire N__43367;
    wire N__43366;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43352;
    wire N__43349;
    wire N__43346;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43331;
    wire N__43328;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43298;
    wire N__43295;
    wire N__43294;
    wire N__43291;
    wire N__43288;
    wire N__43285;
    wire N__43280;
    wire N__43277;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43262;
    wire N__43259;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43244;
    wire N__43241;
    wire N__43240;
    wire N__43237;
    wire N__43234;
    wire N__43231;
    wire N__43226;
    wire N__43223;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43213;
    wire N__43208;
    wire N__43205;
    wire N__43202;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43187;
    wire N__43184;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43169;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43148;
    wire N__43145;
    wire N__43142;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43127;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43115;
    wire N__43112;
    wire N__43109;
    wire N__43106;
    wire N__43103;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43091;
    wire N__43090;
    wire N__43087;
    wire N__43084;
    wire N__43083;
    wire N__43080;
    wire N__43077;
    wire N__43074;
    wire N__43067;
    wire N__43064;
    wire N__43061;
    wire N__43058;
    wire N__43057;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43033;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42995;
    wire N__42992;
    wire N__42989;
    wire N__42986;
    wire N__42983;
    wire N__42980;
    wire N__42977;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42935;
    wire N__42932;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42911;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42854;
    wire N__42851;
    wire N__42848;
    wire N__42845;
    wire N__42842;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42794;
    wire N__42791;
    wire N__42788;
    wire N__42785;
    wire N__42782;
    wire N__42779;
    wire N__42776;
    wire N__42773;
    wire N__42770;
    wire N__42767;
    wire N__42764;
    wire N__42761;
    wire N__42758;
    wire N__42757;
    wire N__42754;
    wire N__42753;
    wire N__42750;
    wire N__42749;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42737;
    wire N__42734;
    wire N__42731;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42715;
    wire N__42710;
    wire N__42707;
    wire N__42704;
    wire N__42701;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42671;
    wire N__42668;
    wire N__42665;
    wire N__42662;
    wire N__42659;
    wire N__42656;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42644;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42626;
    wire N__42623;
    wire N__42620;
    wire N__42617;
    wire N__42614;
    wire N__42611;
    wire N__42608;
    wire N__42605;
    wire N__42602;
    wire N__42599;
    wire N__42596;
    wire N__42593;
    wire N__42590;
    wire N__42587;
    wire N__42584;
    wire N__42581;
    wire N__42578;
    wire N__42575;
    wire N__42572;
    wire N__42571;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42556;
    wire N__42553;
    wire N__42548;
    wire N__42547;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42530;
    wire N__42527;
    wire N__42524;
    wire N__42521;
    wire N__42518;
    wire N__42515;
    wire N__42514;
    wire N__42511;
    wire N__42510;
    wire N__42507;
    wire N__42502;
    wire N__42497;
    wire N__42494;
    wire N__42491;
    wire N__42488;
    wire N__42485;
    wire N__42482;
    wire N__42479;
    wire N__42476;
    wire N__42475;
    wire N__42474;
    wire N__42473;
    wire N__42472;
    wire N__42471;
    wire N__42470;
    wire N__42469;
    wire N__42468;
    wire N__42467;
    wire N__42466;
    wire N__42465;
    wire N__42462;
    wire N__42461;
    wire N__42460;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42452;
    wire N__42451;
    wire N__42448;
    wire N__42447;
    wire N__42446;
    wire N__42445;
    wire N__42444;
    wire N__42443;
    wire N__42442;
    wire N__42441;
    wire N__42440;
    wire N__42439;
    wire N__42438;
    wire N__42437;
    wire N__42434;
    wire N__42433;
    wire N__42432;
    wire N__42431;
    wire N__42428;
    wire N__42425;
    wire N__42424;
    wire N__42423;
    wire N__42422;
    wire N__42421;
    wire N__42420;
    wire N__42417;
    wire N__42416;
    wire N__42413;
    wire N__42412;
    wire N__42411;
    wire N__42408;
    wire N__42407;
    wire N__42404;
    wire N__42403;
    wire N__42400;
    wire N__42399;
    wire N__42398;
    wire N__42397;
    wire N__42396;
    wire N__42395;
    wire N__42394;
    wire N__42393;
    wire N__42392;
    wire N__42391;
    wire N__42390;
    wire N__42389;
    wire N__42388;
    wire N__42387;
    wire N__42384;
    wire N__42373;
    wire N__42370;
    wire N__42359;
    wire N__42342;
    wire N__42339;
    wire N__42328;
    wire N__42327;
    wire N__42326;
    wire N__42325;
    wire N__42324;
    wire N__42323;
    wire N__42322;
    wire N__42321;
    wire N__42320;
    wire N__42319;
    wire N__42318;
    wire N__42315;
    wire N__42314;
    wire N__42311;
    wire N__42310;
    wire N__42307;
    wire N__42306;
    wire N__42305;
    wire N__42304;
    wire N__42303;
    wire N__42302;
    wire N__42301;
    wire N__42300;
    wire N__42299;
    wire N__42298;
    wire N__42297;
    wire N__42296;
    wire N__42291;
    wire N__42274;
    wire N__42265;
    wire N__42262;
    wire N__42261;
    wire N__42258;
    wire N__42257;
    wire N__42254;
    wire N__42253;
    wire N__42250;
    wire N__42249;
    wire N__42248;
    wire N__42247;
    wire N__42246;
    wire N__42245;
    wire N__42244;
    wire N__42243;
    wire N__42242;
    wire N__42241;
    wire N__42238;
    wire N__42237;
    wire N__42234;
    wire N__42233;
    wire N__42230;
    wire N__42229;
    wire N__42226;
    wire N__42225;
    wire N__42222;
    wire N__42221;
    wire N__42218;
    wire N__42217;
    wire N__42214;
    wire N__42213;
    wire N__42208;
    wire N__42205;
    wire N__42200;
    wire N__42195;
    wire N__42188;
    wire N__42185;
    wire N__42184;
    wire N__42183;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42170;
    wire N__42167;
    wire N__42166;
    wire N__42165;
    wire N__42164;
    wire N__42163;
    wire N__42162;
    wire N__42161;
    wire N__42160;
    wire N__42145;
    wire N__42144;
    wire N__42143;
    wire N__42140;
    wire N__42139;
    wire N__42136;
    wire N__42135;
    wire N__42132;
    wire N__42131;
    wire N__42128;
    wire N__42127;
    wire N__42124;
    wire N__42123;
    wire N__42120;
    wire N__42119;
    wire N__42116;
    wire N__42115;
    wire N__42112;
    wire N__42111;
    wire N__42108;
    wire N__42107;
    wire N__42104;
    wire N__42103;
    wire N__42096;
    wire N__42079;
    wire N__42070;
    wire N__42061;
    wire N__42044;
    wire N__42031;
    wire N__42028;
    wire N__42019;
    wire N__42010;
    wire N__42003;
    wire N__42000;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41962;
    wire N__41945;
    wire N__41932;
    wire N__41919;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41885;
    wire N__41882;
    wire N__41879;
    wire N__41878;
    wire N__41875;
    wire N__41874;
    wire N__41867;
    wire N__41864;
    wire N__41863;
    wire N__41862;
    wire N__41861;
    wire N__41860;
    wire N__41859;
    wire N__41858;
    wire N__41857;
    wire N__41856;
    wire N__41855;
    wire N__41854;
    wire N__41853;
    wire N__41852;
    wire N__41849;
    wire N__41848;
    wire N__41847;
    wire N__41846;
    wire N__41845;
    wire N__41844;
    wire N__41843;
    wire N__41840;
    wire N__41827;
    wire N__41816;
    wire N__41813;
    wire N__41808;
    wire N__41807;
    wire N__41806;
    wire N__41805;
    wire N__41804;
    wire N__41803;
    wire N__41802;
    wire N__41793;
    wire N__41786;
    wire N__41781;
    wire N__41778;
    wire N__41767;
    wire N__41760;
    wire N__41753;
    wire N__41750;
    wire N__41749;
    wire N__41748;
    wire N__41745;
    wire N__41742;
    wire N__41739;
    wire N__41732;
    wire N__41729;
    wire N__41728;
    wire N__41727;
    wire N__41724;
    wire N__41721;
    wire N__41718;
    wire N__41711;
    wire N__41708;
    wire N__41705;
    wire N__41702;
    wire N__41699;
    wire N__41698;
    wire N__41695;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41678;
    wire N__41677;
    wire N__41676;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41660;
    wire N__41657;
    wire N__41654;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41646;
    wire N__41641;
    wire N__41638;
    wire N__41633;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41623;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41613;
    wire N__41606;
    wire N__41603;
    wire N__41602;
    wire N__41599;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41572;
    wire N__41569;
    wire N__41566;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41556;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41533;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41516;
    wire N__41515;
    wire N__41512;
    wire N__41509;
    wire N__41508;
    wire N__41503;
    wire N__41500;
    wire N__41495;
    wire N__41492;
    wire N__41491;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41474;
    wire N__41471;
    wire N__41468;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41460;
    wire N__41457;
    wire N__41454;
    wire N__41451;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41429;
    wire N__41426;
    wire N__41425;
    wire N__41424;
    wire N__41421;
    wire N__41416;
    wire N__41411;
    wire N__41408;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41384;
    wire N__41381;
    wire N__41380;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41363;
    wire N__41362;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41352;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41340;
    wire N__41333;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41325;
    wire N__41322;
    wire N__41319;
    wire N__41316;
    wire N__41309;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41292;
    wire N__41285;
    wire N__41284;
    wire N__41283;
    wire N__41280;
    wire N__41277;
    wire N__41276;
    wire N__41273;
    wire N__41270;
    wire N__41267;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41237;
    wire N__41230;
    wire N__41225;
    wire N__41222;
    wire N__41219;
    wire N__41216;
    wire N__41213;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41203;
    wire N__41200;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41183;
    wire N__41182;
    wire N__41181;
    wire N__41176;
    wire N__41173;
    wire N__41168;
    wire N__41167;
    wire N__41164;
    wire N__41161;
    wire N__41160;
    wire N__41157;
    wire N__41154;
    wire N__41151;
    wire N__41144;
    wire N__41141;
    wire N__41140;
    wire N__41137;
    wire N__41134;
    wire N__41131;
    wire N__41126;
    wire N__41123;
    wire N__41122;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41107;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41095;
    wire N__41094;
    wire N__41091;
    wire N__41088;
    wire N__41087;
    wire N__41084;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41061;
    wire N__41058;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41036;
    wire N__41035;
    wire N__41030;
    wire N__41027;
    wire N__41024;
    wire N__41023;
    wire N__41020;
    wire N__41017;
    wire N__41016;
    wire N__41011;
    wire N__41008;
    wire N__41007;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40991;
    wire N__40990;
    wire N__40987;
    wire N__40986;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40966;
    wire N__40961;
    wire N__40960;
    wire N__40959;
    wire N__40956;
    wire N__40953;
    wire N__40950;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40931;
    wire N__40930;
    wire N__40927;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40908;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40894;
    wire N__40889;
    wire N__40888;
    wire N__40887;
    wire N__40884;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40868;
    wire N__40865;
    wire N__40864;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40844;
    wire N__40841;
    wire N__40838;
    wire N__40835;
    wire N__40832;
    wire N__40829;
    wire N__40828;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40813;
    wire N__40808;
    wire N__40805;
    wire N__40804;
    wire N__40803;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40787;
    wire N__40784;
    wire N__40783;
    wire N__40778;
    wire N__40777;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40763;
    wire N__40760;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40748;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40733;
    wire N__40730;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40718;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40693;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40678;
    wire N__40673;
    wire N__40670;
    wire N__40667;
    wire N__40664;
    wire N__40663;
    wire N__40662;
    wire N__40659;
    wire N__40656;
    wire N__40653;
    wire N__40648;
    wire N__40643;
    wire N__40640;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40625;
    wire N__40622;
    wire N__40621;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40606;
    wire N__40601;
    wire N__40598;
    wire N__40597;
    wire N__40596;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40580;
    wire N__40577;
    wire N__40576;
    wire N__40575;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40559;
    wire N__40556;
    wire N__40555;
    wire N__40552;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40537;
    wire N__40532;
    wire N__40529;
    wire N__40528;
    wire N__40525;
    wire N__40524;
    wire N__40521;
    wire N__40518;
    wire N__40515;
    wire N__40510;
    wire N__40505;
    wire N__40502;
    wire N__40501;
    wire N__40498;
    wire N__40495;
    wire N__40494;
    wire N__40489;
    wire N__40486;
    wire N__40483;
    wire N__40478;
    wire N__40475;
    wire N__40474;
    wire N__40471;
    wire N__40468;
    wire N__40467;
    wire N__40462;
    wire N__40459;
    wire N__40456;
    wire N__40451;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40441;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40431;
    wire N__40426;
    wire N__40421;
    wire N__40418;
    wire N__40415;
    wire N__40414;
    wire N__40411;
    wire N__40408;
    wire N__40407;
    wire N__40404;
    wire N__40401;
    wire N__40398;
    wire N__40395;
    wire N__40392;
    wire N__40385;
    wire N__40382;
    wire N__40379;
    wire N__40378;
    wire N__40377;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40363;
    wire N__40358;
    wire N__40355;
    wire N__40354;
    wire N__40353;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40337;
    wire N__40334;
    wire N__40333;
    wire N__40330;
    wire N__40327;
    wire N__40322;
    wire N__40321;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40307;
    wire N__40304;
    wire N__40303;
    wire N__40300;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40290;
    wire N__40285;
    wire N__40280;
    wire N__40279;
    wire N__40278;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40247;
    wire N__40244;
    wire N__40235;
    wire N__40232;
    wire N__40231;
    wire N__40230;
    wire N__40225;
    wire N__40222;
    wire N__40219;
    wire N__40214;
    wire N__40213;
    wire N__40212;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40196;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40172;
    wire N__40169;
    wire N__40168;
    wire N__40165;
    wire N__40162;
    wire N__40161;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40145;
    wire N__40144;
    wire N__40141;
    wire N__40140;
    wire N__40139;
    wire N__40136;
    wire N__40133;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40119;
    wire N__40116;
    wire N__40111;
    wire N__40108;
    wire N__40103;
    wire N__40100;
    wire N__40099;
    wire N__40096;
    wire N__40093;
    wire N__40092;
    wire N__40087;
    wire N__40084;
    wire N__40081;
    wire N__40076;
    wire N__40075;
    wire N__40074;
    wire N__40071;
    wire N__40070;
    wire N__40067;
    wire N__40064;
    wire N__40061;
    wire N__40058;
    wire N__40055;
    wire N__40052;
    wire N__40049;
    wire N__40044;
    wire N__40041;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40025;
    wire N__40024;
    wire N__40023;
    wire N__40020;
    wire N__40017;
    wire N__40014;
    wire N__40009;
    wire N__40004;
    wire N__40003;
    wire N__40002;
    wire N__40001;
    wire N__39998;
    wire N__39995;
    wire N__39992;
    wire N__39989;
    wire N__39986;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39972;
    wire N__39967;
    wire N__39962;
    wire N__39959;
    wire N__39956;
    wire N__39953;
    wire N__39952;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39942;
    wire N__39937;
    wire N__39932;
    wire N__39929;
    wire N__39928;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39920;
    wire N__39917;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39895;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39874;
    wire N__39873;
    wire N__39870;
    wire N__39865;
    wire N__39860;
    wire N__39857;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39847;
    wire N__39842;
    wire N__39839;
    wire N__39838;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39823;
    wire N__39820;
    wire N__39817;
    wire N__39812;
    wire N__39809;
    wire N__39808;
    wire N__39803;
    wire N__39800;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39789;
    wire N__39784;
    wire N__39781;
    wire N__39778;
    wire N__39773;
    wire N__39772;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39764;
    wire N__39761;
    wire N__39758;
    wire N__39755;
    wire N__39750;
    wire N__39743;
    wire N__39740;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39732;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39716;
    wire N__39715;
    wire N__39712;
    wire N__39711;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39699;
    wire N__39696;
    wire N__39691;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39679;
    wire N__39674;
    wire N__39671;
    wire N__39670;
    wire N__39669;
    wire N__39666;
    wire N__39665;
    wire N__39660;
    wire N__39655;
    wire N__39650;
    wire N__39649;
    wire N__39648;
    wire N__39641;
    wire N__39638;
    wire N__39635;
    wire N__39634;
    wire N__39633;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39594;
    wire N__39593;
    wire N__39588;
    wire N__39583;
    wire N__39580;
    wire N__39575;
    wire N__39574;
    wire N__39571;
    wire N__39570;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39547;
    wire N__39542;
    wire N__39539;
    wire N__39538;
    wire N__39537;
    wire N__39536;
    wire N__39535;
    wire N__39534;
    wire N__39525;
    wire N__39524;
    wire N__39523;
    wire N__39522;
    wire N__39521;
    wire N__39520;
    wire N__39519;
    wire N__39518;
    wire N__39517;
    wire N__39516;
    wire N__39515;
    wire N__39514;
    wire N__39513;
    wire N__39512;
    wire N__39511;
    wire N__39510;
    wire N__39509;
    wire N__39508;
    wire N__39507;
    wire N__39506;
    wire N__39505;
    wire N__39504;
    wire N__39503;
    wire N__39502;
    wire N__39501;
    wire N__39496;
    wire N__39493;
    wire N__39484;
    wire N__39475;
    wire N__39466;
    wire N__39457;
    wire N__39448;
    wire N__39439;
    wire N__39436;
    wire N__39431;
    wire N__39418;
    wire N__39415;
    wire N__39412;
    wire N__39407;
    wire N__39406;
    wire N__39405;
    wire N__39402;
    wire N__39397;
    wire N__39396;
    wire N__39391;
    wire N__39388;
    wire N__39385;
    wire N__39380;
    wire N__39379;
    wire N__39376;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39338;
    wire N__39335;
    wire N__39334;
    wire N__39331;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39315;
    wire N__39308;
    wire N__39307;
    wire N__39304;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39288;
    wire N__39281;
    wire N__39280;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39259;
    wire N__39254;
    wire N__39253;
    wire N__39252;
    wire N__39251;
    wire N__39248;
    wire N__39243;
    wire N__39240;
    wire N__39235;
    wire N__39230;
    wire N__39229;
    wire N__39228;
    wire N__39227;
    wire N__39220;
    wire N__39219;
    wire N__39216;
    wire N__39215;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39195;
    wire N__39188;
    wire N__39183;
    wire N__39180;
    wire N__39173;
    wire N__39172;
    wire N__39169;
    wire N__39168;
    wire N__39167;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39152;
    wire N__39143;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39116;
    wire N__39113;
    wire N__39110;
    wire N__39107;
    wire N__39106;
    wire N__39103;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39086;
    wire N__39083;
    wire N__39080;
    wire N__39079;
    wire N__39076;
    wire N__39075;
    wire N__39072;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39056;
    wire N__39053;
    wire N__39050;
    wire N__39047;
    wire N__39044;
    wire N__39041;
    wire N__39038;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38990;
    wire N__38987;
    wire N__38984;
    wire N__38981;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38973;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38941;
    wire N__38940;
    wire N__38937;
    wire N__38932;
    wire N__38927;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38915;
    wire N__38912;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38904;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38892;
    wire N__38889;
    wire N__38882;
    wire N__38879;
    wire N__38876;
    wire N__38873;
    wire N__38872;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38846;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38834;
    wire N__38831;
    wire N__38828;
    wire N__38827;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38804;
    wire N__38801;
    wire N__38798;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38735;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38717;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38702;
    wire N__38699;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38674;
    wire N__38671;
    wire N__38666;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38651;
    wire N__38650;
    wire N__38647;
    wire N__38642;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38627;
    wire N__38626;
    wire N__38621;
    wire N__38618;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38582;
    wire N__38579;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38558;
    wire N__38557;
    wire N__38554;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38543;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38519;
    wire N__38516;
    wire N__38515;
    wire N__38512;
    wire N__38509;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38473;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38456;
    wire N__38455;
    wire N__38452;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38429;
    wire N__38426;
    wire N__38423;
    wire N__38420;
    wire N__38417;
    wire N__38414;
    wire N__38411;
    wire N__38408;
    wire N__38405;
    wire N__38404;
    wire N__38403;
    wire N__38400;
    wire N__38395;
    wire N__38390;
    wire N__38389;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38377;
    wire N__38372;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38354;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38321;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38267;
    wire N__38264;
    wire N__38261;
    wire N__38260;
    wire N__38259;
    wire N__38256;
    wire N__38251;
    wire N__38246;
    wire N__38243;
    wire N__38242;
    wire N__38241;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38225;
    wire N__38222;
    wire N__38219;
    wire N__38216;
    wire N__38213;
    wire N__38210;
    wire N__38209;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38197;
    wire N__38192;
    wire N__38189;
    wire N__38186;
    wire N__38183;
    wire N__38180;
    wire N__38177;
    wire N__38174;
    wire N__38171;
    wire N__38168;
    wire N__38165;
    wire N__38162;
    wire N__38159;
    wire N__38156;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38132;
    wire N__38131;
    wire N__38130;
    wire N__38129;
    wire N__38128;
    wire N__38127;
    wire N__38126;
    wire N__38125;
    wire N__38124;
    wire N__38123;
    wire N__38122;
    wire N__38121;
    wire N__38120;
    wire N__38119;
    wire N__38118;
    wire N__38117;
    wire N__38108;
    wire N__38099;
    wire N__38098;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38094;
    wire N__38093;
    wire N__38092;
    wire N__38091;
    wire N__38090;
    wire N__38089;
    wire N__38088;
    wire N__38087;
    wire N__38086;
    wire N__38085;
    wire N__38076;
    wire N__38067;
    wire N__38062;
    wire N__38053;
    wire N__38048;
    wire N__38039;
    wire N__38030;
    wire N__38025;
    wire N__38014;
    wire N__38009;
    wire N__38006;
    wire N__38003;
    wire N__38002;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37991;
    wire N__37988;
    wire N__37983;
    wire N__37980;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37958;
    wire N__37955;
    wire N__37952;
    wire N__37949;
    wire N__37946;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37880;
    wire N__37877;
    wire N__37874;
    wire N__37871;
    wire N__37868;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37838;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37805;
    wire N__37802;
    wire N__37799;
    wire N__37796;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37778;
    wire N__37775;
    wire N__37772;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37666;
    wire N__37665;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37653;
    wire N__37646;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37591;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37502;
    wire N__37499;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37484;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37436;
    wire N__37435;
    wire N__37434;
    wire N__37433;
    wire N__37432;
    wire N__37431;
    wire N__37430;
    wire N__37429;
    wire N__37428;
    wire N__37427;
    wire N__37426;
    wire N__37425;
    wire N__37424;
    wire N__37423;
    wire N__37422;
    wire N__37421;
    wire N__37420;
    wire N__37419;
    wire N__37418;
    wire N__37417;
    wire N__37416;
    wire N__37415;
    wire N__37414;
    wire N__37413;
    wire N__37410;
    wire N__37409;
    wire N__37408;
    wire N__37407;
    wire N__37406;
    wire N__37405;
    wire N__37404;
    wire N__37403;
    wire N__37402;
    wire N__37393;
    wire N__37384;
    wire N__37377;
    wire N__37368;
    wire N__37359;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37337;
    wire N__37328;
    wire N__37323;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37299;
    wire N__37296;
    wire N__37289;
    wire N__37286;
    wire N__37285;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37273;
    wire N__37270;
    wire N__37269;
    wire N__37268;
    wire N__37267;
    wire N__37264;
    wire N__37261;
    wire N__37254;
    wire N__37247;
    wire N__37244;
    wire N__37243;
    wire N__37242;
    wire N__37239;
    wire N__37236;
    wire N__37233;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37066;
    wire N__37063;
    wire N__37060;
    wire N__37055;
    wire N__37052;
    wire N__37051;
    wire N__37050;
    wire N__37049;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36994;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36911;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36878;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36866;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36833;
    wire N__36830;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36806;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36754;
    wire N__36751;
    wire N__36748;
    wire N__36745;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36730;
    wire N__36727;
    wire N__36724;
    wire N__36721;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36700;
    wire N__36697;
    wire N__36694;
    wire N__36691;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36661;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36640;
    wire N__36637;
    wire N__36634;
    wire N__36631;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36610;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36598;
    wire N__36597;
    wire N__36594;
    wire N__36589;
    wire N__36584;
    wire N__36581;
    wire N__36580;
    wire N__36579;
    wire N__36574;
    wire N__36571;
    wire N__36568;
    wire N__36563;
    wire N__36560;
    wire N__36559;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36538;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36511;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36499;
    wire N__36494;
    wire N__36491;
    wire N__36490;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36478;
    wire N__36473;
    wire N__36470;
    wire N__36469;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36457;
    wire N__36452;
    wire N__36449;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36419;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36406;
    wire N__36405;
    wire N__36402;
    wire N__36397;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36337;
    wire N__36336;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36304;
    wire N__36301;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36284;
    wire N__36281;
    wire N__36280;
    wire N__36277;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36260;
    wire N__36259;
    wire N__36256;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36203;
    wire N__36200;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36176;
    wire N__36173;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36101;
    wire N__36098;
    wire N__36095;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35918;
    wire N__35915;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35881;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35873;
    wire N__35872;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35850;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35825;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35813;
    wire N__35812;
    wire N__35811;
    wire N__35808;
    wire N__35805;
    wire N__35804;
    wire N__35801;
    wire N__35796;
    wire N__35793;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35764;
    wire N__35763;
    wire N__35760;
    wire N__35757;
    wire N__35754;
    wire N__35749;
    wire N__35744;
    wire N__35743;
    wire N__35740;
    wire N__35739;
    wire N__35736;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35724;
    wire N__35721;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35709;
    wire N__35702;
    wire N__35701;
    wire N__35700;
    wire N__35699;
    wire N__35696;
    wire N__35689;
    wire N__35686;
    wire N__35681;
    wire N__35680;
    wire N__35679;
    wire N__35676;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35651;
    wire N__35650;
    wire N__35647;
    wire N__35646;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35636;
    wire N__35633;
    wire N__35628;
    wire N__35625;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35608;
    wire N__35607;
    wire N__35604;
    wire N__35599;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35569;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35554;
    wire N__35549;
    wire N__35548;
    wire N__35543;
    wire N__35540;
    wire N__35539;
    wire N__35534;
    wire N__35531;
    wire N__35530;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35518;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35495;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35473;
    wire N__35472;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35461;
    wire N__35458;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35441;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35427;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35404;
    wire N__35403;
    wire N__35402;
    wire N__35401;
    wire N__35400;
    wire N__35399;
    wire N__35398;
    wire N__35397;
    wire N__35396;
    wire N__35395;
    wire N__35392;
    wire N__35391;
    wire N__35388;
    wire N__35385;
    wire N__35384;
    wire N__35383;
    wire N__35382;
    wire N__35381;
    wire N__35380;
    wire N__35377;
    wire N__35376;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35358;
    wire N__35355;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35343;
    wire N__35340;
    wire N__35339;
    wire N__35338;
    wire N__35337;
    wire N__35336;
    wire N__35335;
    wire N__35334;
    wire N__35333;
    wire N__35332;
    wire N__35331;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35320;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35302;
    wire N__35293;
    wire N__35292;
    wire N__35289;
    wire N__35282;
    wire N__35279;
    wire N__35274;
    wire N__35261;
    wire N__35254;
    wire N__35253;
    wire N__35240;
    wire N__35239;
    wire N__35238;
    wire N__35237;
    wire N__35236;
    wire N__35235;
    wire N__35234;
    wire N__35233;
    wire N__35232;
    wire N__35231;
    wire N__35228;
    wire N__35221;
    wire N__35218;
    wire N__35217;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35178;
    wire N__35177;
    wire N__35176;
    wire N__35175;
    wire N__35174;
    wire N__35171;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35151;
    wire N__35142;
    wire N__35129;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35121;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35098;
    wire N__35093;
    wire N__35092;
    wire N__35089;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35066;
    wire N__35065;
    wire N__35062;
    wire N__35059;
    wire N__35058;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35016;
    wire N__35011;
    wire N__35006;
    wire N__35003;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34962;
    wire N__34961;
    wire N__34960;
    wire N__34955;
    wire N__34948;
    wire N__34943;
    wire N__34942;
    wire N__34941;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34904;
    wire N__34903;
    wire N__34902;
    wire N__34899;
    wire N__34894;
    wire N__34889;
    wire N__34888;
    wire N__34885;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34841;
    wire N__34838;
    wire N__34837;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34820;
    wire N__34819;
    wire N__34818;
    wire N__34811;
    wire N__34806;
    wire N__34803;
    wire N__34796;
    wire N__34793;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34768;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34745;
    wire N__34744;
    wire N__34743;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34724;
    wire N__34721;
    wire N__34716;
    wire N__34713;
    wire N__34706;
    wire N__34705;
    wire N__34704;
    wire N__34703;
    wire N__34702;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34698;
    wire N__34697;
    wire N__34696;
    wire N__34695;
    wire N__34694;
    wire N__34693;
    wire N__34690;
    wire N__34689;
    wire N__34688;
    wire N__34687;
    wire N__34686;
    wire N__34685;
    wire N__34684;
    wire N__34683;
    wire N__34682;
    wire N__34681;
    wire N__34680;
    wire N__34679;
    wire N__34678;
    wire N__34677;
    wire N__34676;
    wire N__34675;
    wire N__34674;
    wire N__34673;
    wire N__34672;
    wire N__34669;
    wire N__34668;
    wire N__34667;
    wire N__34666;
    wire N__34665;
    wire N__34664;
    wire N__34663;
    wire N__34662;
    wire N__34651;
    wire N__34642;
    wire N__34629;
    wire N__34626;
    wire N__34625;
    wire N__34624;
    wire N__34623;
    wire N__34622;
    wire N__34617;
    wire N__34616;
    wire N__34615;
    wire N__34614;
    wire N__34613;
    wire N__34612;
    wire N__34611;
    wire N__34610;
    wire N__34609;
    wire N__34608;
    wire N__34607;
    wire N__34606;
    wire N__34605;
    wire N__34604;
    wire N__34603;
    wire N__34602;
    wire N__34599;
    wire N__34598;
    wire N__34597;
    wire N__34596;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34592;
    wire N__34591;
    wire N__34590;
    wire N__34589;
    wire N__34588;
    wire N__34587;
    wire N__34586;
    wire N__34579;
    wire N__34578;
    wire N__34577;
    wire N__34576;
    wire N__34575;
    wire N__34562;
    wire N__34551;
    wire N__34538;
    wire N__34533;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34521;
    wire N__34516;
    wire N__34515;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34511;
    wire N__34508;
    wire N__34501;
    wire N__34496;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34484;
    wire N__34483;
    wire N__34482;
    wire N__34481;
    wire N__34480;
    wire N__34477;
    wire N__34476;
    wire N__34473;
    wire N__34472;
    wire N__34471;
    wire N__34470;
    wire N__34469;
    wire N__34468;
    wire N__34457;
    wire N__34454;
    wire N__34441;
    wire N__34430;
    wire N__34427;
    wire N__34424;
    wire N__34415;
    wire N__34406;
    wire N__34403;
    wire N__34396;
    wire N__34393;
    wire N__34382;
    wire N__34377;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34359;
    wire N__34354;
    wire N__34349;
    wire N__34346;
    wire N__34335;
    wire N__34326;
    wire N__34317;
    wire N__34312;
    wire N__34301;
    wire N__34298;
    wire N__34291;
    wire N__34274;
    wire N__34273;
    wire N__34270;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34258;
    wire N__34255;
    wire N__34254;
    wire N__34253;
    wire N__34252;
    wire N__34251;
    wire N__34250;
    wire N__34249;
    wire N__34248;
    wire N__34247;
    wire N__34246;
    wire N__34245;
    wire N__34244;
    wire N__34243;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34207;
    wire N__34206;
    wire N__34205;
    wire N__34204;
    wire N__34203;
    wire N__34202;
    wire N__34201;
    wire N__34200;
    wire N__34199;
    wire N__34196;
    wire N__34193;
    wire N__34192;
    wire N__34191;
    wire N__34190;
    wire N__34189;
    wire N__34186;
    wire N__34185;
    wire N__34184;
    wire N__34183;
    wire N__34182;
    wire N__34181;
    wire N__34180;
    wire N__34179;
    wire N__34178;
    wire N__34177;
    wire N__34176;
    wire N__34175;
    wire N__34170;
    wire N__34167;
    wire N__34166;
    wire N__34165;
    wire N__34164;
    wire N__34163;
    wire N__34156;
    wire N__34155;
    wire N__34152;
    wire N__34145;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34095;
    wire N__34086;
    wire N__34081;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34058;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34039;
    wire N__34032;
    wire N__34025;
    wire N__34018;
    wire N__34009;
    wire N__34006;
    wire N__34001;
    wire N__33998;
    wire N__33995;
    wire N__33986;
    wire N__33983;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33887;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33839;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33825;
    wire N__33820;
    wire N__33817;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33692;
    wire N__33691;
    wire N__33690;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33641;
    wire N__33638;
    wire N__33637;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33622;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33584;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33572;
    wire N__33571;
    wire N__33566;
    wire N__33565;
    wire N__33564;
    wire N__33561;
    wire N__33556;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33524;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33481;
    wire N__33478;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33432;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33416;
    wire N__33413;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33405;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33389;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33343;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33328;
    wire N__33323;
    wire N__33320;
    wire N__33319;
    wire N__33318;
    wire N__33315;
    wire N__33312;
    wire N__33309;
    wire N__33304;
    wire N__33299;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33236;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33188;
    wire N__33187;
    wire N__33186;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33056;
    wire N__33053;
    wire N__33052;
    wire N__33049;
    wire N__33046;
    wire N__33041;
    wire N__33038;
    wire N__33035;
    wire N__33032;
    wire N__33029;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33007;
    wire N__33006;
    wire N__33003;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32987;
    wire N__32984;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32933;
    wire N__32930;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32922;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32900;
    wire N__32891;
    wire N__32888;
    wire N__32887;
    wire N__32884;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32867;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32852;
    wire N__32849;
    wire N__32848;
    wire N__32843;
    wire N__32842;
    wire N__32839;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32809;
    wire N__32806;
    wire N__32805;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32787;
    wire N__32784;
    wire N__32777;
    wire N__32774;
    wire N__32773;
    wire N__32770;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32731;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32713;
    wire N__32708;
    wire N__32707;
    wire N__32704;
    wire N__32701;
    wire N__32700;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32682;
    wire N__32679;
    wire N__32672;
    wire N__32671;
    wire N__32666;
    wire N__32663;
    wire N__32662;
    wire N__32659;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32642;
    wire N__32639;
    wire N__32638;
    wire N__32635;
    wire N__32634;
    wire N__32631;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32584;
    wire N__32581;
    wire N__32580;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32564;
    wire N__32563;
    wire N__32562;
    wire N__32559;
    wire N__32554;
    wire N__32549;
    wire N__32548;
    wire N__32545;
    wire N__32540;
    wire N__32537;
    wire N__32536;
    wire N__32533;
    wire N__32530;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32516;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32503;
    wire N__32500;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32483;
    wire N__32480;
    wire N__32479;
    wire N__32476;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32459;
    wire N__32456;
    wire N__32455;
    wire N__32452;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32428;
    wire N__32425;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32398;
    wire N__32397;
    wire N__32396;
    wire N__32395;
    wire N__32394;
    wire N__32393;
    wire N__32392;
    wire N__32391;
    wire N__32390;
    wire N__32389;
    wire N__32388;
    wire N__32387;
    wire N__32386;
    wire N__32385;
    wire N__32384;
    wire N__32383;
    wire N__32382;
    wire N__32381;
    wire N__32380;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32369;
    wire N__32368;
    wire N__32367;
    wire N__32366;
    wire N__32365;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32353;
    wire N__32352;
    wire N__32351;
    wire N__32350;
    wire N__32343;
    wire N__32332;
    wire N__32329;
    wire N__32328;
    wire N__32327;
    wire N__32326;
    wire N__32323;
    wire N__32320;
    wire N__32309;
    wire N__32306;
    wire N__32299;
    wire N__32292;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32259;
    wire N__32254;
    wire N__32249;
    wire N__32246;
    wire N__32241;
    wire N__32238;
    wire N__32225;
    wire N__32224;
    wire N__32223;
    wire N__32220;
    wire N__32219;
    wire N__32216;
    wire N__32215;
    wire N__32214;
    wire N__32213;
    wire N__32212;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32204;
    wire N__32203;
    wire N__32202;
    wire N__32201;
    wire N__32200;
    wire N__32199;
    wire N__32198;
    wire N__32197;
    wire N__32194;
    wire N__32193;
    wire N__32192;
    wire N__32189;
    wire N__32188;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32158;
    wire N__32157;
    wire N__32156;
    wire N__32155;
    wire N__32154;
    wire N__32153;
    wire N__32142;
    wire N__32135;
    wire N__32134;
    wire N__32133;
    wire N__32132;
    wire N__32131;
    wire N__32130;
    wire N__32127;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32103;
    wire N__32096;
    wire N__32089;
    wire N__32084;
    wire N__32073;
    wire N__32068;
    wire N__32065;
    wire N__32056;
    wire N__32053;
    wire N__32048;
    wire N__32045;
    wire N__32042;
    wire N__32033;
    wire N__32032;
    wire N__32031;
    wire N__32030;
    wire N__32029;
    wire N__32028;
    wire N__32027;
    wire N__32026;
    wire N__32025;
    wire N__32024;
    wire N__32023;
    wire N__32022;
    wire N__32021;
    wire N__32020;
    wire N__32019;
    wire N__32018;
    wire N__32017;
    wire N__32016;
    wire N__32015;
    wire N__32014;
    wire N__32013;
    wire N__32010;
    wire N__32009;
    wire N__32006;
    wire N__32005;
    wire N__32004;
    wire N__32003;
    wire N__32000;
    wire N__31993;
    wire N__31992;
    wire N__31981;
    wire N__31970;
    wire N__31959;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31949;
    wire N__31948;
    wire N__31947;
    wire N__31946;
    wire N__31945;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31922;
    wire N__31919;
    wire N__31912;
    wire N__31901;
    wire N__31894;
    wire N__31887;
    wire N__31884;
    wire N__31879;
    wire N__31868;
    wire N__31865;
    wire N__31864;
    wire N__31861;
    wire N__31858;
    wire N__31857;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31847;
    wire N__31844;
    wire N__31843;
    wire N__31838;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31798;
    wire N__31797;
    wire N__31796;
    wire N__31795;
    wire N__31794;
    wire N__31791;
    wire N__31790;
    wire N__31787;
    wire N__31786;
    wire N__31783;
    wire N__31782;
    wire N__31779;
    wire N__31778;
    wire N__31761;
    wire N__31760;
    wire N__31759;
    wire N__31758;
    wire N__31757;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31745;
    wire N__31742;
    wire N__31741;
    wire N__31738;
    wire N__31737;
    wire N__31734;
    wire N__31733;
    wire N__31730;
    wire N__31727;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31691;
    wire N__31688;
    wire N__31685;
    wire N__31682;
    wire N__31681;
    wire N__31680;
    wire N__31677;
    wire N__31672;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31654;
    wire N__31651;
    wire N__31650;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31490;
    wire N__31489;
    wire N__31486;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31469;
    wire N__31466;
    wire N__31465;
    wire N__31462;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31445;
    wire N__31442;
    wire N__31441;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31418;
    wire N__31415;
    wire N__31414;
    wire N__31411;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31357;
    wire N__31354;
    wire N__31351;
    wire N__31348;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31304;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31280;
    wire N__31277;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31235;
    wire N__31232;
    wire N__31229;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31202;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31172;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31147;
    wire N__31144;
    wire N__31141;
    wire N__31138;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31121;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31009;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30994;
    wire N__30991;
    wire N__30988;
    wire N__30985;
    wire N__30980;
    wire N__30977;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30955;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30931;
    wire N__30930;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30907;
    wire N__30906;
    wire N__30905;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30880;
    wire N__30879;
    wire N__30878;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30860;
    wire N__30857;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30784;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30706;
    wire N__30703;
    wire N__30702;
    wire N__30699;
    wire N__30694;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30682;
    wire N__30677;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30662;
    wire N__30659;
    wire N__30658;
    wire N__30657;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30641;
    wire N__30638;
    wire N__30637;
    wire N__30636;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30620;
    wire N__30617;
    wire N__30616;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30592;
    wire N__30589;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30566;
    wire N__30563;
    wire N__30562;
    wire N__30559;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30542;
    wire N__30539;
    wire N__30538;
    wire N__30535;
    wire N__30534;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30518;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30497;
    wire N__30496;
    wire N__30493;
    wire N__30492;
    wire N__30489;
    wire N__30484;
    wire N__30479;
    wire N__30476;
    wire N__30475;
    wire N__30474;
    wire N__30471;
    wire N__30466;
    wire N__30461;
    wire N__30458;
    wire N__30457;
    wire N__30456;
    wire N__30453;
    wire N__30448;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30434;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30403;
    wire N__30400;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30390;
    wire N__30383;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30368;
    wire N__30365;
    wire N__30360;
    wire N__30357;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30337;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30316;
    wire N__30313;
    wire N__30312;
    wire N__30309;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30274;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30242;
    wire N__30239;
    wire N__30238;
    wire N__30235;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30200;
    wire N__30197;
    wire N__30196;
    wire N__30195;
    wire N__30192;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30171;
    wire N__30164;
    wire N__30161;
    wire N__30160;
    wire N__30155;
    wire N__30152;
    wire N__30151;
    wire N__30148;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30131;
    wire N__30130;
    wire N__30127;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30113;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30095;
    wire N__30094;
    wire N__30091;
    wire N__30090;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30054;
    wire N__30051;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30025;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30005;
    wire N__30004;
    wire N__30001;
    wire N__30000;
    wire N__29997;
    wire N__29994;
    wire N__29991;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29977;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29966;
    wire N__29965;
    wire N__29962;
    wire N__29957;
    wire N__29952;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29935;
    wire N__29932;
    wire N__29931;
    wire N__29928;
    wire N__29925;
    wire N__29922;
    wire N__29915;
    wire N__29914;
    wire N__29911;
    wire N__29910;
    wire N__29909;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29885;
    wire N__29880;
    wire N__29875;
    wire N__29872;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29839;
    wire N__29836;
    wire N__29835;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29789;
    wire N__29784;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29767;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29756;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29729;
    wire N__29726;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29690;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29561;
    wire N__29558;
    wire N__29555;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29446;
    wire N__29445;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29433;
    wire N__29428;
    wire N__29425;
    wire N__29420;
    wire N__29417;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29405;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29393;
    wire N__29392;
    wire N__29389;
    wire N__29386;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29326;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29289;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29277;
    wire N__29270;
    wire N__29267;
    wire N__29266;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29243;
    wire N__29240;
    wire N__29237;
    wire N__29236;
    wire N__29235;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29223;
    wire N__29216;
    wire N__29213;
    wire N__29210;
    wire N__29209;
    wire N__29206;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29189;
    wire N__29188;
    wire N__29185;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29163;
    wire N__29156;
    wire N__29153;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29141;
    wire N__29140;
    wire N__29139;
    wire N__29136;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29101;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29075;
    wire N__29074;
    wire N__29073;
    wire N__29068;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29058;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29005;
    wire N__29004;
    wire N__29003;
    wire N__29000;
    wire N__28995;
    wire N__28992;
    wire N__28985;
    wire N__28982;
    wire N__28981;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28955;
    wire N__28952;
    wire N__28949;
    wire N__28948;
    wire N__28947;
    wire N__28944;
    wire N__28939;
    wire N__28938;
    wire N__28933;
    wire N__28930;
    wire N__28925;
    wire N__28924;
    wire N__28919;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28898;
    wire N__28895;
    wire N__28894;
    wire N__28893;
    wire N__28890;
    wire N__28885;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28868;
    wire N__28867;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28852;
    wire N__28851;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28836;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28815;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28803;
    wire N__28796;
    wire N__28793;
    wire N__28792;
    wire N__28791;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28779;
    wire N__28776;
    wire N__28769;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28744;
    wire N__28743;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28731;
    wire N__28728;
    wire N__28721;
    wire N__28720;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28706;
    wire N__28703;
    wire N__28702;
    wire N__28701;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28676;
    wire N__28675;
    wire N__28674;
    wire N__28673;
    wire N__28670;
    wire N__28665;
    wire N__28662;
    wire N__28655;
    wire N__28654;
    wire N__28651;
    wire N__28650;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28638;
    wire N__28631;
    wire N__28630;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28607;
    wire N__28606;
    wire N__28605;
    wire N__28604;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28562;
    wire N__28559;
    wire N__28558;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28547;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28493;
    wire N__28490;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28455;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28443;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28422;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28381;
    wire N__28380;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28368;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28340;
    wire N__28337;
    wire N__28336;
    wire N__28335;
    wire N__28334;
    wire N__28331;
    wire N__28324;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28297;
    wire N__28294;
    wire N__28293;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28272;
    wire N__28269;
    wire N__28264;
    wire N__28261;
    wire N__28258;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28234;
    wire N__28233;
    wire N__28230;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28209;
    wire N__28206;
    wire N__28205;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28187;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28179;
    wire N__28176;
    wire N__28171;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28150;
    wire N__28147;
    wire N__28144;
    wire N__28139;
    wire N__28136;
    wire N__28135;
    wire N__28134;
    wire N__28131;
    wire N__28126;
    wire N__28123;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28053;
    wire N__28052;
    wire N__28049;
    wire N__28044;
    wire N__28043;
    wire N__28040;
    wire N__28035;
    wire N__28032;
    wire N__28027;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28012;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27983;
    wire N__27980;
    wire N__27975;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27939;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27931;
    wire N__27926;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27866;
    wire N__27863;
    wire N__27862;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27854;
    wire N__27851;
    wire N__27846;
    wire N__27843;
    wire N__27838;
    wire N__27837;
    wire N__27832;
    wire N__27829;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27817;
    wire N__27814;
    wire N__27813;
    wire N__27810;
    wire N__27809;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27783;
    wire N__27780;
    wire N__27775;
    wire N__27772;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27748;
    wire N__27745;
    wire N__27744;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27709;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27694;
    wire N__27693;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27685;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27658;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27634;
    wire N__27631;
    wire N__27630;
    wire N__27629;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27560;
    wire N__27559;
    wire N__27556;
    wire N__27551;
    wire N__27546;
    wire N__27543;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27529;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27518;
    wire N__27515;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27488;
    wire N__27485;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27443;
    wire N__27440;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27423;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27409;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27388;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27370;
    wire N__27369;
    wire N__27366;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27330;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27260;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27242;
    wire N__27241;
    wire N__27240;
    wire N__27237;
    wire N__27232;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27202;
    wire N__27201;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27157;
    wire N__27154;
    wire N__27153;
    wire N__27150;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27132;
    wire N__27131;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27084;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27072;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27049;
    wire N__27048;
    wire N__27045;
    wire N__27040;
    wire N__27035;
    wire N__27034;
    wire N__27033;
    wire N__27030;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26989;
    wire N__26988;
    wire N__26987;
    wire N__26984;
    wire N__26979;
    wire N__26976;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26945;
    wire N__26942;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26879;
    wire N__26876;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26865;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26853;
    wire N__26850;
    wire N__26843;
    wire N__26842;
    wire N__26839;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26827;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26804;
    wire N__26803;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26791;
    wire N__26788;
    wire N__26787;
    wire N__26786;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26772;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26758;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26744;
    wire N__26743;
    wire N__26740;
    wire N__26737;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26729;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26714;
    wire N__26705;
    wire N__26704;
    wire N__26703;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26658;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26642;
    wire N__26639;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26625;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26602;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26587;
    wire N__26582;
    wire N__26579;
    wire N__26578;
    wire N__26577;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26561;
    wire N__26558;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26522;
    wire N__26519;
    wire N__26518;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26503;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26491;
    wire N__26490;
    wire N__26487;
    wire N__26484;
    wire N__26483;
    wire N__26480;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26444;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26432;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26424;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26412;
    wire N__26407;
    wire N__26402;
    wire N__26399;
    wire N__26398;
    wire N__26393;
    wire N__26392;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26378;
    wire N__26375;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26367;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26351;
    wire N__26348;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26334;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26308;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26298;
    wire N__26293;
    wire N__26288;
    wire N__26285;
    wire N__26284;
    wire N__26283;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26267;
    wire N__26264;
    wire N__26263;
    wire N__26262;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26246;
    wire N__26243;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26235;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26219;
    wire N__26216;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26208;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26192;
    wire N__26189;
    wire N__26188;
    wire N__26183;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26168;
    wire N__26167;
    wire N__26162;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26147;
    wire N__26144;
    wire N__26143;
    wire N__26138;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26123;
    wire N__26120;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26106;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26090;
    wire N__26087;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26065;
    wire N__26060;
    wire N__26057;
    wire N__26056;
    wire N__26051;
    wire N__26050;
    wire N__26047;
    wire N__26044;
    wire N__26041;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26022;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26006;
    wire N__26003;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25995;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25979;
    wire N__25976;
    wire N__25975;
    wire N__25974;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25948;
    wire N__25947;
    wire N__25946;
    wire N__25945;
    wire N__25944;
    wire N__25943;
    wire N__25942;
    wire N__25941;
    wire N__25940;
    wire N__25939;
    wire N__25938;
    wire N__25937;
    wire N__25936;
    wire N__25935;
    wire N__25934;
    wire N__25933;
    wire N__25932;
    wire N__25931;
    wire N__25930;
    wire N__25929;
    wire N__25928;
    wire N__25927;
    wire N__25926;
    wire N__25925;
    wire N__25924;
    wire N__25923;
    wire N__25922;
    wire N__25921;
    wire N__25920;
    wire N__25911;
    wire N__25902;
    wire N__25893;
    wire N__25888;
    wire N__25879;
    wire N__25870;
    wire N__25861;
    wire N__25852;
    wire N__25845;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25818;
    wire N__25813;
    wire N__25810;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25795;
    wire N__25792;
    wire N__25787;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25776;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25760;
    wire N__25757;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25749;
    wire N__25744;
    wire N__25741;
    wire N__25736;
    wire N__25733;
    wire N__25732;
    wire N__25727;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25712;
    wire N__25709;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25684;
    wire N__25679;
    wire N__25676;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25668;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25652;
    wire N__25649;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25641;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25491;
    wire N__25488;
    wire N__25487;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24994;
    wire N__24993;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24981;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24964;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24952;
    wire N__24951;
    wire N__24948;
    wire N__24943;
    wire N__24938;
    wire N__24935;
    wire N__24934;
    wire N__24933;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24917;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24892;
    wire N__24891;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24875;
    wire N__24872;
    wire N__24871;
    wire N__24870;
    wire N__24865;
    wire N__24862;
    wire N__24859;
    wire N__24854;
    wire N__24853;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24826;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24814;
    wire N__24809;
    wire N__24806;
    wire N__24805;
    wire N__24804;
    wire N__24803;
    wire N__24802;
    wire N__24801;
    wire N__24800;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24775;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24718;
    wire N__24715;
    wire N__24714;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24702;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24664;
    wire N__24661;
    wire N__24660;
    wire N__24657;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24628;
    wire N__24627;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24611;
    wire N__24608;
    wire N__24607;
    wire N__24602;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24580;
    wire N__24575;
    wire N__24572;
    wire N__24569;
    wire N__24568;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24514;
    wire N__24513;
    wire N__24506;
    wire N__24503;
    wire N__24502;
    wire N__24501;
    wire N__24498;
    wire N__24491;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24476;
    wire N__24475;
    wire N__24474;
    wire N__24467;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24433;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24415;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24376;
    wire N__24371;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24356;
    wire N__24353;
    wire N__24352;
    wire N__24347;
    wire N__24344;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24322;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24310;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24283;
    wire N__24278;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24263;
    wire N__24260;
    wire N__24259;
    wire N__24254;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24226;
    wire N__24225;
    wire N__24224;
    wire N__24221;
    wire N__24214;
    wire N__24209;
    wire N__24206;
    wire N__24205;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24190;
    wire N__24189;
    wire N__24188;
    wire N__24183;
    wire N__24178;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24131;
    wire N__24130;
    wire N__24127;
    wire N__24122;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24098;
    wire N__24097;
    wire N__24096;
    wire N__24095;
    wire N__24094;
    wire N__24093;
    wire N__24092;
    wire N__24091;
    wire N__24090;
    wire N__24089;
    wire N__24088;
    wire N__24087;
    wire N__24078;
    wire N__24071;
    wire N__24062;
    wire N__24053;
    wire N__24052;
    wire N__24051;
    wire N__24050;
    wire N__24049;
    wire N__24048;
    wire N__24047;
    wire N__24046;
    wire N__24045;
    wire N__24044;
    wire N__24043;
    wire N__24042;
    wire N__24041;
    wire N__24040;
    wire N__24039;
    wire N__24038;
    wire N__24037;
    wire N__24034;
    wire N__24027;
    wire N__24020;
    wire N__24011;
    wire N__24002;
    wire N__23993;
    wire N__23990;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23886;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23870;
    wire N__23867;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23852;
    wire N__23849;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23813;
    wire N__23810;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23795;
    wire N__23792;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23767;
    wire N__23766;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23743;
    wire N__23738;
    wire N__23737;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23723;
    wire N__23720;
    wire N__23719;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23705;
    wire N__23702;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23645;
    wire N__23642;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23627;
    wire N__23624;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23533;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23518;
    wire N__23513;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23308;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23296;
    wire N__23291;
    wire N__23288;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23276;
    wire N__23273;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23191;
    wire N__23190;
    wire N__23189;
    wire N__23188;
    wire N__23187;
    wire N__23184;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23169;
    wire N__23168;
    wire N__23167;
    wire N__23166;
    wire N__23155;
    wire N__23152;
    wire N__23147;
    wire N__23144;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23110;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23060;
    wire N__23057;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23042;
    wire N__23039;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23009;
    wire N__23006;
    wire N__23005;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22993;
    wire N__22990;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22957;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22921;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22909;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22861;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22838;
    wire N__22835;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22816;
    wire N__22813;
    wire N__22810;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22753;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22711;
    wire N__22708;
    wire N__22707;
    wire N__22704;
    wire N__22703;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22675;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22647;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22564;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22513;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22463;
    wire N__22462;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22408;
    wire N__22407;
    wire N__22406;
    wire N__22405;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22377;
    wire N__22376;
    wire N__22373;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22296;
    wire N__22295;
    wire N__22294;
    wire N__22293;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22281;
    wire N__22280;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22266;
    wire N__22261;
    wire N__22258;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22236;
    wire N__22233;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22117;
    wire N__22116;
    wire N__22115;
    wire N__22114;
    wire N__22111;
    wire N__22110;
    wire N__22109;
    wire N__22100;
    wire N__22099;
    wire N__22098;
    wire N__22097;
    wire N__22094;
    wire N__22089;
    wire N__22086;
    wire N__22079;
    wire N__22074;
    wire N__22069;
    wire N__22066;
    wire N__22061;
    wire N__22060;
    wire N__22059;
    wire N__22058;
    wire N__22057;
    wire N__22054;
    wire N__22053;
    wire N__22050;
    wire N__22049;
    wire N__22048;
    wire N__22045;
    wire N__22044;
    wire N__22041;
    wire N__22040;
    wire N__22037;
    wire N__22032;
    wire N__22029;
    wire N__22020;
    wire N__22013;
    wire N__22012;
    wire N__22011;
    wire N__22010;
    wire N__22009;
    wire N__22008;
    wire N__21999;
    wire N__21998;
    wire N__21997;
    wire N__21996;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21985;
    wire N__21984;
    wire N__21979;
    wire N__21972;
    wire N__21969;
    wire N__21968;
    wire N__21951;
    wire N__21936;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21924;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21886;
    wire N__21885;
    wire N__21884;
    wire N__21883;
    wire N__21882;
    wire N__21881;
    wire N__21872;
    wire N__21865;
    wire N__21864;
    wire N__21863;
    wire N__21862;
    wire N__21857;
    wire N__21850;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21803;
    wire N__21800;
    wire N__21799;
    wire N__21796;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21781;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21757;
    wire N__21754;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21586;
    wire N__21583;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21550;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21535;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21518;
    wire N__21517;
    wire N__21516;
    wire N__21515;
    wire N__21514;
    wire N__21513;
    wire N__21512;
    wire N__21503;
    wire N__21494;
    wire N__21489;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21473;
    wire N__21472;
    wire N__21471;
    wire N__21470;
    wire N__21467;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21379;
    wire N__21376;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21283;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21268;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21238;
    wire N__21235;
    wire N__21234;
    wire N__21231;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21220;
    wire N__21219;
    wire N__21218;
    wire N__21215;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21205;
    wire N__21204;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21196;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21178;
    wire N__21165;
    wire N__21158;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21128;
    wire N__21125;
    wire N__21124;
    wire N__21121;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21104;
    wire N__21101;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21082;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21062;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21044;
    wire N__21041;
    wire N__21040;
    wire N__21037;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20770;
    wire N__20769;
    wire N__20766;
    wire N__20761;
    wire N__20756;
    wire N__20753;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20695;
    wire N__20692;
    wire N__20689;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20584;
    wire N__20583;
    wire N__20580;
    wire N__20575;
    wire N__20572;
    wire N__20567;
    wire N__20566;
    wire N__20565;
    wire N__20560;
    wire N__20557;
    wire N__20552;
    wire N__20549;
    wire N__20548;
    wire N__20545;
    wire N__20544;
    wire N__20541;
    wire N__20538;
    wire N__20533;
    wire N__20530;
    wire N__20525;
    wire N__20522;
    wire N__20521;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20494;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20474;
    wire N__20471;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20456;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20444;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20404;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20386;
    wire N__20381;
    wire N__20380;
    wire N__20379;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20362;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20287;
    wire N__20286;
    wire N__20281;
    wire N__20278;
    wire N__20273;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20161;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20128;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20089;
    wire N__20086;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19882;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19801;
    wire N__19796;
    wire N__19793;
    wire N__19792;
    wire N__19791;
    wire N__19790;
    wire N__19789;
    wire N__19788;
    wire N__19787;
    wire N__19784;
    wire N__19777;
    wire N__19770;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19396;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire bfn_1_9_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_1_10_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire bfn_1_13_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire bfn_1_14_0_;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire bfn_1_15_0_;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10_cascade_ ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_1_19_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_1_20_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire bfn_1_21_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire N_42_i_i;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire pwm_duty_input_7;
    wire pwm_duty_input_5;
    wire pwm_duty_input_6;
    wire pwm_duty_input_8;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_3;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ;
    wire pwm_duty_input_4;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \current_shift_inst.PI_CTRL.N_140 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_145 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire bfn_2_14_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ;
    wire bfn_2_15_0_;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0 ;
    wire bfn_2_16_0_;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire bfn_2_17_0_;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791 ;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire bfn_2_18_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire un7_start_stop_0_a2;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto9_2_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9 ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \current_shift_inst.PI_CTRL.N_144 ;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31 ;
    wire \current_shift_inst.PI_CTRL.N_146 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61 ;
    wire \pwm_generator_inst.threshold_0 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_3_15_0_;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_3_16_0_;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671 ;
    wire \pwm_generator_inst.threshold_9 ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61 ;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.N_16 ;
    wire N_19_1;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1 ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_53 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_71 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ;
    wire \current_shift_inst.PI_CTRL.un1_enablelt3_0 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_164 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_5_15_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_5_16_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_5_17_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_5_18_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_7_9_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_7_10_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire bfn_7_11_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_7_12_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_7_13_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_7_14_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_7_15_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_72_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13_cascade_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12_cascade_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26_cascade_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.un1_start_g ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire bfn_8_16_0_;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire bfn_8_17_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire bfn_8_18_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_30 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_30 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire s4_phy_c;
    wire bfn_9_4_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_9_5_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_9_6_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_9_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_204_i ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_9_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_9_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_9_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_9_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_203_i ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27_cascade_;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire elapsed_time_ns_1_RNI6HPBB_0_28_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_ ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.state_RNIG7JFZ0Z_2_cascade_ ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire s3_phy_c;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire il_max_comp1_c;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire elapsed_time_ns_1_RNIU7OBB_0_11_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire elapsed_time_ns_1_RNILK91B_0_9_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire elapsed_time_ns_1_RNIVAQBB_0_30_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire elapsed_time_ns_1_RNI0CQBB_0_31_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire elapsed_time_ns_1_RNI6GOBB_0_19_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire elapsed_time_ns_1_RNI5FOBB_0_18_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire elapsed_time_ns_1_RNIU8PBB_0_20_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ;
    wire bfn_10_14_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_8 ;
    wire bfn_10_15_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ;
    wire bfn_10_16_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ;
    wire bfn_10_17_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_31 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ;
    wire il_min_comp1_c;
    wire il_max_comp1_D1;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire elapsed_time_ns_1_RNI1CPBB_0_23_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df30 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire bfn_11_9_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire bfn_11_10_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_11_11_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire bfn_11_12_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_11_13_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_11_14_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire bfn_11_15_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.N_74 ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire il_max_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire il_min_comp1_D1;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire elapsed_time_ns_1_RNI1BOBB_0_14_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire bfn_12_11_0_;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire bfn_12_12_0_;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.control_input_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_12_13_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_12_14_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ;
    wire \phase_controller_inst1.N_55_cascade_ ;
    wire state_ns_i_a2_1;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ;
    wire \phase_controller_inst2.state_RNIG7JFZ0Z_2 ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire T23_c;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire T45_c;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.N_1326_i ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.control_input_axb_9 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ;
    wire \phase_controller_inst1.N_55 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire start_stop_c;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst1.N_54 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire T12_c;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_19 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire \current_shift_inst.timer_s1.N_167_i ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire s1_phy_c;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire delay_hc_input_c_g;
    wire bfn_14_5_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire bfn_14_6_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_14_7_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_14_8_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire bfn_14_9_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire bfn_14_10_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_14_11_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_14_12_0_;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \pll_inst.red_c_i ;
    wire il_max_comp1_D2;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire bfn_14_19_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_14_20_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_14_21_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_14_22_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_14_24_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_14_25_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire bfn_14_26_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire bfn_15_13_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire bfn_15_14_0_;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire bfn_15_15_0_;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire bfn_15_16_0_;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.N_168_i ;
    wire bfn_15_17_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_15_18_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_15_19_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_15_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt30 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire bfn_16_8_0_;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_16_9_0_;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire bfn_16_10_0_;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_16_11_0_;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_202_i ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire \phase_controller_inst1.hc_time_passed ;
    wire state_3;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire T01_c;
    wire \phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire elapsed_time_ns_1_RNI14DN9_0_23_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire elapsed_time_ns_1_RNI03DN9_0_22_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire bfn_16_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire bfn_16_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_16_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_16_23_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_201_i ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_11 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_17_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_17_16_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire bfn_17_17_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire bfn_17_18_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_17_19_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_17_20_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_17_21_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire elapsed_time_ns_1_RNI7ADN9_0_29_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire bfn_18_7_0_;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_18_8_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire bfn_18_9_0_;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire bfn_18_10_0_;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire bfn_18_11_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire bfn_18_12_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire bfn_18_13_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire bfn_18_14_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.N_167_i_g ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire elapsed_time_ns_1_RNI46CN9_0_17_cascade_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire elapsed_time_ns_1_RNI13CN9_0_14_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire elapsed_time_ns_1_RNI25DN9_0_24_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire elapsed_time_ns_1_RNI57CN9_0_18_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire \phase_controller_inst2.stoper_hc.un1_start_g ;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__28088),
            .RESETB(N__36362),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__44988),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__44981),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__21997,N__21990,N__21995,N__21989,N__21996,N__21988,N__21998,N__21985,N__21991,N__21984,N__21992,N__21986,N__21993,N__21987,N__21994}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__44987,N__44984,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__44982,N__44986,N__44983,N__44985}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__44925),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__44873),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .ADDSUBBOT(),
            .A({dangling_wire_74,N__22010,N__22012,N__22008,N__22011,N__22009,N__20549,N__20565,N__20286,N__20588,N__20273,N__20498,N__20525,N__20443,N__20455,N__20474}),
            .C({dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90}),
            .B({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__44879,N__44876,dangling_wire_98,dangling_wire_99,dangling_wire_100,N__44874,N__44878,N__44875,N__44877}),
            .OHOLDTOP(),
            .O({dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__50430),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__50432),
            .DIN(N__50431),
            .DOUT(N__50430),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__50432),
            .PADOUT(N__50431),
            .PADIN(N__50430),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__50421),
            .DIN(N__50420),
            .DOUT(N__50419),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__50421),
            .PADOUT(N__50420),
            .PADIN(N__50419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__39143),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__50412),
            .DIN(N__50411),
            .DOUT(N__50410),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__50412),
            .PADOUT(N__50411),
            .PADIN(N__50410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__50403),
            .DIN(N__50402),
            .DOUT(N__50401),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__50403),
            .PADOUT(N__50402),
            .PADIN(N__50401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__50394),
            .DIN(N__50393),
            .DOUT(N__50392),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__50394),
            .PADOUT(N__50393),
            .PADIN(N__50392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33596),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__50385),
            .DIN(N__50384),
            .DOUT(N__50383),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__50385),
            .PADOUT(N__50384),
            .PADIN(N__50383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22196),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__50376),
            .DIN(N__50375),
            .DOUT(N__50374),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__50376),
            .PADOUT(N__50375),
            .PADIN(N__50374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__50367),
            .DIN(N__50366),
            .DOUT(N__50365),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__50367),
            .PADOUT(N__50366),
            .PADIN(N__50365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35837),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__50358),
            .DIN(N__50357),
            .DOUT(N__50356),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__50358),
            .PADOUT(N__50357),
            .PADIN(N__50356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35510),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__50349),
            .DIN(N__50348),
            .DOUT(N__50347),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__50349),
            .PADOUT(N__50348),
            .PADIN(N__50347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__50340),
            .DIN(N__50339),
            .DOUT(N__50338),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__50340),
            .PADOUT(N__50339),
            .PADIN(N__50338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__50331),
            .DIN(N__50330),
            .DOUT(N__50329),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__50331),
            .PADOUT(N__50330),
            .PADIN(N__50329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25445),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__50322),
            .DIN(N__50321),
            .DOUT(N__50320),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__50322),
            .PADOUT(N__50321),
            .PADIN(N__50320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__50313),
            .DIN(N__50312),
            .DOUT(N__50311),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__50313),
            .PADOUT(N__50312),
            .PADIN(N__50311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28109),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__50304),
            .DIN(N__50303),
            .DOUT(N__50302),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__50304),
            .PADOUT(N__50303),
            .PADIN(N__50302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33551),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__50295),
            .DIN(N__50294),
            .DOUT(N__50293),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__50295),
            .PADOUT(N__50294),
            .PADIN(N__50293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__50286),
            .DIN(N__50285),
            .DOUT(N__50284),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__50286),
            .PADOUT(N__50285),
            .PADIN(N__50284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11929 (
            .O(N__50267),
            .I(N__50264));
    LocalMux I__11928 (
            .O(N__50264),
            .I(N__50261));
    Span4Mux_v I__11927 (
            .O(N__50261),
            .I(N__50255));
    InMux I__11926 (
            .O(N__50260),
            .I(N__50252));
    InMux I__11925 (
            .O(N__50259),
            .I(N__50249));
    InMux I__11924 (
            .O(N__50258),
            .I(N__50246));
    Odrv4 I__11923 (
            .O(N__50255),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    LocalMux I__11922 (
            .O(N__50252),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    LocalMux I__11921 (
            .O(N__50249),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    LocalMux I__11920 (
            .O(N__50246),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__11919 (
            .O(N__50237),
            .I(N__50232));
    InMux I__11918 (
            .O(N__50236),
            .I(N__50229));
    InMux I__11917 (
            .O(N__50235),
            .I(N__50226));
    LocalMux I__11916 (
            .O(N__50232),
            .I(N__50223));
    LocalMux I__11915 (
            .O(N__50229),
            .I(N__50220));
    LocalMux I__11914 (
            .O(N__50226),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__11913 (
            .O(N__50223),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__11912 (
            .O(N__50220),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    CascadeMux I__11911 (
            .O(N__50213),
            .I(N__50209));
    CascadeMux I__11910 (
            .O(N__50212),
            .I(N__50206));
    InMux I__11909 (
            .O(N__50209),
            .I(N__50201));
    InMux I__11908 (
            .O(N__50206),
            .I(N__50201));
    LocalMux I__11907 (
            .O(N__50201),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ));
    InMux I__11906 (
            .O(N__50198),
            .I(N__50194));
    InMux I__11905 (
            .O(N__50197),
            .I(N__50190));
    LocalMux I__11904 (
            .O(N__50194),
            .I(N__50187));
    InMux I__11903 (
            .O(N__50193),
            .I(N__50184));
    LocalMux I__11902 (
            .O(N__50190),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    Odrv12 I__11901 (
            .O(N__50187),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    LocalMux I__11900 (
            .O(N__50184),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    InMux I__11899 (
            .O(N__50177),
            .I(N__50174));
    LocalMux I__11898 (
            .O(N__50174),
            .I(N__50169));
    InMux I__11897 (
            .O(N__50173),
            .I(N__50166));
    InMux I__11896 (
            .O(N__50172),
            .I(N__50163));
    Span4Mux_v I__11895 (
            .O(N__50169),
            .I(N__50157));
    LocalMux I__11894 (
            .O(N__50166),
            .I(N__50157));
    LocalMux I__11893 (
            .O(N__50163),
            .I(N__50154));
    InMux I__11892 (
            .O(N__50162),
            .I(N__50151));
    Odrv4 I__11891 (
            .O(N__50157),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__11890 (
            .O(N__50154),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__11889 (
            .O(N__50151),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__11888 (
            .O(N__50144),
            .I(N__50138));
    InMux I__11887 (
            .O(N__50143),
            .I(N__50138));
    LocalMux I__11886 (
            .O(N__50138),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ));
    InMux I__11885 (
            .O(N__50135),
            .I(N__50129));
    InMux I__11884 (
            .O(N__50134),
            .I(N__50126));
    InMux I__11883 (
            .O(N__50133),
            .I(N__50121));
    InMux I__11882 (
            .O(N__50132),
            .I(N__50121));
    LocalMux I__11881 (
            .O(N__50129),
            .I(N__50118));
    LocalMux I__11880 (
            .O(N__50126),
            .I(N__50115));
    LocalMux I__11879 (
            .O(N__50121),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__11878 (
            .O(N__50118),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__11877 (
            .O(N__50115),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    CascadeMux I__11876 (
            .O(N__50108),
            .I(N__50105));
    InMux I__11875 (
            .O(N__50105),
            .I(N__50102));
    LocalMux I__11874 (
            .O(N__50102),
            .I(N__50095));
    InMux I__11873 (
            .O(N__50101),
            .I(N__50092));
    InMux I__11872 (
            .O(N__50100),
            .I(N__50089));
    InMux I__11871 (
            .O(N__50099),
            .I(N__50084));
    InMux I__11870 (
            .O(N__50098),
            .I(N__50084));
    Span4Mux_v I__11869 (
            .O(N__50095),
            .I(N__50079));
    LocalMux I__11868 (
            .O(N__50092),
            .I(N__50079));
    LocalMux I__11867 (
            .O(N__50089),
            .I(N__50074));
    LocalMux I__11866 (
            .O(N__50084),
            .I(N__50074));
    Span4Mux_h I__11865 (
            .O(N__50079),
            .I(N__50071));
    Odrv12 I__11864 (
            .O(N__50074),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__11863 (
            .O(N__50071),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    CEMux I__11862 (
            .O(N__50066),
            .I(N__50063));
    LocalMux I__11861 (
            .O(N__50063),
            .I(N__50059));
    CEMux I__11860 (
            .O(N__50062),
            .I(N__50056));
    Span4Mux_v I__11859 (
            .O(N__50059),
            .I(N__50042));
    LocalMux I__11858 (
            .O(N__50056),
            .I(N__50042));
    InMux I__11857 (
            .O(N__50055),
            .I(N__50035));
    InMux I__11856 (
            .O(N__50054),
            .I(N__50035));
    InMux I__11855 (
            .O(N__50053),
            .I(N__50035));
    InMux I__11854 (
            .O(N__50052),
            .I(N__50028));
    InMux I__11853 (
            .O(N__50051),
            .I(N__50018));
    InMux I__11852 (
            .O(N__50050),
            .I(N__50018));
    InMux I__11851 (
            .O(N__50049),
            .I(N__50018));
    InMux I__11850 (
            .O(N__50048),
            .I(N__50018));
    CEMux I__11849 (
            .O(N__50047),
            .I(N__50015));
    Span4Mux_h I__11848 (
            .O(N__50042),
            .I(N__50010));
    LocalMux I__11847 (
            .O(N__50035),
            .I(N__50010));
    CEMux I__11846 (
            .O(N__50034),
            .I(N__50007));
    CEMux I__11845 (
            .O(N__50033),
            .I(N__50002));
    CEMux I__11844 (
            .O(N__50032),
            .I(N__49995));
    CEMux I__11843 (
            .O(N__50031),
            .I(N__49991));
    LocalMux I__11842 (
            .O(N__50028),
            .I(N__49987));
    CEMux I__11841 (
            .O(N__50027),
            .I(N__49984));
    LocalMux I__11840 (
            .O(N__50018),
            .I(N__49970));
    LocalMux I__11839 (
            .O(N__50015),
            .I(N__49970));
    Span4Mux_v I__11838 (
            .O(N__50010),
            .I(N__49965));
    LocalMux I__11837 (
            .O(N__50007),
            .I(N__49965));
    CEMux I__11836 (
            .O(N__50006),
            .I(N__49949));
    CEMux I__11835 (
            .O(N__50005),
            .I(N__49946));
    LocalMux I__11834 (
            .O(N__50002),
            .I(N__49943));
    InMux I__11833 (
            .O(N__50001),
            .I(N__49934));
    InMux I__11832 (
            .O(N__50000),
            .I(N__49934));
    InMux I__11831 (
            .O(N__49999),
            .I(N__49934));
    InMux I__11830 (
            .O(N__49998),
            .I(N__49934));
    LocalMux I__11829 (
            .O(N__49995),
            .I(N__49931));
    CEMux I__11828 (
            .O(N__49994),
            .I(N__49928));
    LocalMux I__11827 (
            .O(N__49991),
            .I(N__49925));
    CEMux I__11826 (
            .O(N__49990),
            .I(N__49922));
    Span4Mux_v I__11825 (
            .O(N__49987),
            .I(N__49917));
    LocalMux I__11824 (
            .O(N__49984),
            .I(N__49917));
    CEMux I__11823 (
            .O(N__49983),
            .I(N__49914));
    CEMux I__11822 (
            .O(N__49982),
            .I(N__49911));
    InMux I__11821 (
            .O(N__49981),
            .I(N__49902));
    InMux I__11820 (
            .O(N__49980),
            .I(N__49902));
    InMux I__11819 (
            .O(N__49979),
            .I(N__49902));
    InMux I__11818 (
            .O(N__49978),
            .I(N__49902));
    InMux I__11817 (
            .O(N__49977),
            .I(N__49895));
    InMux I__11816 (
            .O(N__49976),
            .I(N__49895));
    InMux I__11815 (
            .O(N__49975),
            .I(N__49895));
    Span4Mux_v I__11814 (
            .O(N__49970),
            .I(N__49890));
    Span4Mux_v I__11813 (
            .O(N__49965),
            .I(N__49890));
    InMux I__11812 (
            .O(N__49964),
            .I(N__49881));
    InMux I__11811 (
            .O(N__49963),
            .I(N__49881));
    InMux I__11810 (
            .O(N__49962),
            .I(N__49881));
    InMux I__11809 (
            .O(N__49961),
            .I(N__49881));
    InMux I__11808 (
            .O(N__49960),
            .I(N__49872));
    InMux I__11807 (
            .O(N__49959),
            .I(N__49872));
    InMux I__11806 (
            .O(N__49958),
            .I(N__49872));
    InMux I__11805 (
            .O(N__49957),
            .I(N__49872));
    InMux I__11804 (
            .O(N__49956),
            .I(N__49863));
    InMux I__11803 (
            .O(N__49955),
            .I(N__49863));
    InMux I__11802 (
            .O(N__49954),
            .I(N__49863));
    InMux I__11801 (
            .O(N__49953),
            .I(N__49863));
    CEMux I__11800 (
            .O(N__49952),
            .I(N__49860));
    LocalMux I__11799 (
            .O(N__49949),
            .I(N__49855));
    LocalMux I__11798 (
            .O(N__49946),
            .I(N__49855));
    Span4Mux_h I__11797 (
            .O(N__49943),
            .I(N__49852));
    LocalMux I__11796 (
            .O(N__49934),
            .I(N__49849));
    Span4Mux_h I__11795 (
            .O(N__49931),
            .I(N__49846));
    LocalMux I__11794 (
            .O(N__49928),
            .I(N__49837));
    Span4Mux_h I__11793 (
            .O(N__49925),
            .I(N__49837));
    LocalMux I__11792 (
            .O(N__49922),
            .I(N__49837));
    Span4Mux_h I__11791 (
            .O(N__49917),
            .I(N__49837));
    LocalMux I__11790 (
            .O(N__49914),
            .I(N__49834));
    LocalMux I__11789 (
            .O(N__49911),
            .I(N__49831));
    LocalMux I__11788 (
            .O(N__49902),
            .I(N__49818));
    LocalMux I__11787 (
            .O(N__49895),
            .I(N__49818));
    Span4Mux_h I__11786 (
            .O(N__49890),
            .I(N__49818));
    LocalMux I__11785 (
            .O(N__49881),
            .I(N__49818));
    LocalMux I__11784 (
            .O(N__49872),
            .I(N__49818));
    LocalMux I__11783 (
            .O(N__49863),
            .I(N__49818));
    LocalMux I__11782 (
            .O(N__49860),
            .I(N__49815));
    Span4Mux_h I__11781 (
            .O(N__49855),
            .I(N__49810));
    Span4Mux_h I__11780 (
            .O(N__49852),
            .I(N__49810));
    Span4Mux_h I__11779 (
            .O(N__49849),
            .I(N__49801));
    Span4Mux_h I__11778 (
            .O(N__49846),
            .I(N__49801));
    Span4Mux_h I__11777 (
            .O(N__49837),
            .I(N__49801));
    Span4Mux_h I__11776 (
            .O(N__49834),
            .I(N__49801));
    Span12Mux_h I__11775 (
            .O(N__49831),
            .I(N__49798));
    Span4Mux_v I__11774 (
            .O(N__49818),
            .I(N__49795));
    Span4Mux_h I__11773 (
            .O(N__49815),
            .I(N__49790));
    Span4Mux_v I__11772 (
            .O(N__49810),
            .I(N__49790));
    Span4Mux_v I__11771 (
            .O(N__49801),
            .I(N__49787));
    Odrv12 I__11770 (
            .O(N__49798),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11769 (
            .O(N__49795),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11768 (
            .O(N__49790),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11767 (
            .O(N__49787),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__11766 (
            .O(N__49778),
            .I(N__49774));
    CascadeMux I__11765 (
            .O(N__49777),
            .I(N__49770));
    LocalMux I__11764 (
            .O(N__49774),
            .I(N__49766));
    InMux I__11763 (
            .O(N__49773),
            .I(N__49763));
    InMux I__11762 (
            .O(N__49770),
            .I(N__49760));
    InMux I__11761 (
            .O(N__49769),
            .I(N__49757));
    Span4Mux_h I__11760 (
            .O(N__49766),
            .I(N__49754));
    LocalMux I__11759 (
            .O(N__49763),
            .I(N__49749));
    LocalMux I__11758 (
            .O(N__49760),
            .I(N__49749));
    LocalMux I__11757 (
            .O(N__49757),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__11756 (
            .O(N__49754),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv12 I__11755 (
            .O(N__49749),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__11754 (
            .O(N__49742),
            .I(N__49738));
    InMux I__11753 (
            .O(N__49741),
            .I(N__49735));
    LocalMux I__11752 (
            .O(N__49738),
            .I(N__49731));
    LocalMux I__11751 (
            .O(N__49735),
            .I(N__49728));
    InMux I__11750 (
            .O(N__49734),
            .I(N__49725));
    Span4Mux_h I__11749 (
            .O(N__49731),
            .I(N__49720));
    Span4Mux_v I__11748 (
            .O(N__49728),
            .I(N__49720));
    LocalMux I__11747 (
            .O(N__49725),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    Odrv4 I__11746 (
            .O(N__49720),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__11745 (
            .O(N__49715),
            .I(N__49710));
    InMux I__11744 (
            .O(N__49714),
            .I(N__49706));
    InMux I__11743 (
            .O(N__49713),
            .I(N__49703));
    LocalMux I__11742 (
            .O(N__49710),
            .I(N__49700));
    InMux I__11741 (
            .O(N__49709),
            .I(N__49697));
    LocalMux I__11740 (
            .O(N__49706),
            .I(N__49694));
    LocalMux I__11739 (
            .O(N__49703),
            .I(N__49691));
    Span4Mux_v I__11738 (
            .O(N__49700),
            .I(N__49688));
    LocalMux I__11737 (
            .O(N__49697),
            .I(N__49685));
    Span4Mux_v I__11736 (
            .O(N__49694),
            .I(N__49682));
    Span12Mux_s9_h I__11735 (
            .O(N__49691),
            .I(N__49679));
    Span4Mux_h I__11734 (
            .O(N__49688),
            .I(N__49674));
    Span4Mux_h I__11733 (
            .O(N__49685),
            .I(N__49674));
    Odrv4 I__11732 (
            .O(N__49682),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv12 I__11731 (
            .O(N__49679),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__11730 (
            .O(N__49674),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__11729 (
            .O(N__49667),
            .I(N__49663));
    InMux I__11728 (
            .O(N__49666),
            .I(N__49660));
    LocalMux I__11727 (
            .O(N__49663),
            .I(N__49656));
    LocalMux I__11726 (
            .O(N__49660),
            .I(N__49653));
    InMux I__11725 (
            .O(N__49659),
            .I(N__49650));
    Span4Mux_v I__11724 (
            .O(N__49656),
            .I(N__49645));
    Span4Mux_h I__11723 (
            .O(N__49653),
            .I(N__49645));
    LocalMux I__11722 (
            .O(N__49650),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    Odrv4 I__11721 (
            .O(N__49645),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    InMux I__11720 (
            .O(N__49640),
            .I(N__49632));
    InMux I__11719 (
            .O(N__49639),
            .I(N__49620));
    InMux I__11718 (
            .O(N__49638),
            .I(N__49604));
    InMux I__11717 (
            .O(N__49637),
            .I(N__49604));
    InMux I__11716 (
            .O(N__49636),
            .I(N__49604));
    InMux I__11715 (
            .O(N__49635),
            .I(N__49604));
    LocalMux I__11714 (
            .O(N__49632),
            .I(N__49601));
    InMux I__11713 (
            .O(N__49631),
            .I(N__49594));
    InMux I__11712 (
            .O(N__49630),
            .I(N__49594));
    InMux I__11711 (
            .O(N__49629),
            .I(N__49594));
    InMux I__11710 (
            .O(N__49628),
            .I(N__49556));
    InMux I__11709 (
            .O(N__49627),
            .I(N__49556));
    InMux I__11708 (
            .O(N__49626),
            .I(N__49556));
    InMux I__11707 (
            .O(N__49625),
            .I(N__49556));
    InMux I__11706 (
            .O(N__49624),
            .I(N__49556));
    CascadeMux I__11705 (
            .O(N__49623),
            .I(N__49551));
    LocalMux I__11704 (
            .O(N__49620),
            .I(N__49543));
    InMux I__11703 (
            .O(N__49619),
            .I(N__49538));
    InMux I__11702 (
            .O(N__49618),
            .I(N__49538));
    InMux I__11701 (
            .O(N__49617),
            .I(N__49535));
    InMux I__11700 (
            .O(N__49616),
            .I(N__49527));
    InMux I__11699 (
            .O(N__49615),
            .I(N__49520));
    InMux I__11698 (
            .O(N__49614),
            .I(N__49520));
    InMux I__11697 (
            .O(N__49613),
            .I(N__49520));
    LocalMux I__11696 (
            .O(N__49604),
            .I(N__49517));
    Span4Mux_h I__11695 (
            .O(N__49601),
            .I(N__49512));
    LocalMux I__11694 (
            .O(N__49594),
            .I(N__49512));
    InMux I__11693 (
            .O(N__49593),
            .I(N__49509));
    InMux I__11692 (
            .O(N__49592),
            .I(N__49498));
    InMux I__11691 (
            .O(N__49591),
            .I(N__49498));
    InMux I__11690 (
            .O(N__49590),
            .I(N__49498));
    InMux I__11689 (
            .O(N__49589),
            .I(N__49498));
    InMux I__11688 (
            .O(N__49588),
            .I(N__49498));
    InMux I__11687 (
            .O(N__49587),
            .I(N__49489));
    InMux I__11686 (
            .O(N__49586),
            .I(N__49489));
    InMux I__11685 (
            .O(N__49585),
            .I(N__49489));
    InMux I__11684 (
            .O(N__49584),
            .I(N__49489));
    InMux I__11683 (
            .O(N__49583),
            .I(N__49482));
    InMux I__11682 (
            .O(N__49582),
            .I(N__49482));
    InMux I__11681 (
            .O(N__49581),
            .I(N__49482));
    InMux I__11680 (
            .O(N__49580),
            .I(N__49476));
    CascadeMux I__11679 (
            .O(N__49579),
            .I(N__49473));
    CascadeMux I__11678 (
            .O(N__49578),
            .I(N__49470));
    InMux I__11677 (
            .O(N__49577),
            .I(N__49466));
    InMux I__11676 (
            .O(N__49576),
            .I(N__49459));
    InMux I__11675 (
            .O(N__49575),
            .I(N__49459));
    InMux I__11674 (
            .O(N__49574),
            .I(N__49459));
    InMux I__11673 (
            .O(N__49573),
            .I(N__49447));
    InMux I__11672 (
            .O(N__49572),
            .I(N__49447));
    InMux I__11671 (
            .O(N__49571),
            .I(N__49436));
    InMux I__11670 (
            .O(N__49570),
            .I(N__49436));
    InMux I__11669 (
            .O(N__49569),
            .I(N__49436));
    InMux I__11668 (
            .O(N__49568),
            .I(N__49436));
    InMux I__11667 (
            .O(N__49567),
            .I(N__49436));
    LocalMux I__11666 (
            .O(N__49556),
            .I(N__49433));
    InMux I__11665 (
            .O(N__49555),
            .I(N__49430));
    InMux I__11664 (
            .O(N__49554),
            .I(N__49426));
    InMux I__11663 (
            .O(N__49551),
            .I(N__49415));
    InMux I__11662 (
            .O(N__49550),
            .I(N__49408));
    InMux I__11661 (
            .O(N__49549),
            .I(N__49408));
    InMux I__11660 (
            .O(N__49548),
            .I(N__49408));
    InMux I__11659 (
            .O(N__49547),
            .I(N__49403));
    InMux I__11658 (
            .O(N__49546),
            .I(N__49403));
    Span4Mux_v I__11657 (
            .O(N__49543),
            .I(N__49400));
    LocalMux I__11656 (
            .O(N__49538),
            .I(N__49395));
    LocalMux I__11655 (
            .O(N__49535),
            .I(N__49395));
    InMux I__11654 (
            .O(N__49534),
            .I(N__49392));
    InMux I__11653 (
            .O(N__49533),
            .I(N__49383));
    InMux I__11652 (
            .O(N__49532),
            .I(N__49383));
    InMux I__11651 (
            .O(N__49531),
            .I(N__49383));
    InMux I__11650 (
            .O(N__49530),
            .I(N__49383));
    LocalMux I__11649 (
            .O(N__49527),
            .I(N__49372));
    LocalMux I__11648 (
            .O(N__49520),
            .I(N__49372));
    Span4Mux_v I__11647 (
            .O(N__49517),
            .I(N__49372));
    Span4Mux_v I__11646 (
            .O(N__49512),
            .I(N__49372));
    LocalMux I__11645 (
            .O(N__49509),
            .I(N__49372));
    LocalMux I__11644 (
            .O(N__49498),
            .I(N__49367));
    LocalMux I__11643 (
            .O(N__49489),
            .I(N__49367));
    LocalMux I__11642 (
            .O(N__49482),
            .I(N__49364));
    InMux I__11641 (
            .O(N__49481),
            .I(N__49357));
    InMux I__11640 (
            .O(N__49480),
            .I(N__49357));
    InMux I__11639 (
            .O(N__49479),
            .I(N__49357));
    LocalMux I__11638 (
            .O(N__49476),
            .I(N__49354));
    InMux I__11637 (
            .O(N__49473),
            .I(N__49343));
    InMux I__11636 (
            .O(N__49470),
            .I(N__49343));
    InMux I__11635 (
            .O(N__49469),
            .I(N__49343));
    LocalMux I__11634 (
            .O(N__49466),
            .I(N__49340));
    LocalMux I__11633 (
            .O(N__49459),
            .I(N__49337));
    InMux I__11632 (
            .O(N__49458),
            .I(N__49329));
    InMux I__11631 (
            .O(N__49457),
            .I(N__49329));
    InMux I__11630 (
            .O(N__49456),
            .I(N__49322));
    InMux I__11629 (
            .O(N__49455),
            .I(N__49322));
    InMux I__11628 (
            .O(N__49454),
            .I(N__49322));
    InMux I__11627 (
            .O(N__49453),
            .I(N__49313));
    InMux I__11626 (
            .O(N__49452),
            .I(N__49313));
    LocalMux I__11625 (
            .O(N__49447),
            .I(N__49304));
    LocalMux I__11624 (
            .O(N__49436),
            .I(N__49304));
    Sp12to4 I__11623 (
            .O(N__49433),
            .I(N__49304));
    LocalMux I__11622 (
            .O(N__49430),
            .I(N__49304));
    InMux I__11621 (
            .O(N__49429),
            .I(N__49301));
    LocalMux I__11620 (
            .O(N__49426),
            .I(N__49298));
    InMux I__11619 (
            .O(N__49425),
            .I(N__49295));
    InMux I__11618 (
            .O(N__49424),
            .I(N__49288));
    InMux I__11617 (
            .O(N__49423),
            .I(N__49288));
    InMux I__11616 (
            .O(N__49422),
            .I(N__49288));
    InMux I__11615 (
            .O(N__49421),
            .I(N__49281));
    InMux I__11614 (
            .O(N__49420),
            .I(N__49281));
    InMux I__11613 (
            .O(N__49419),
            .I(N__49281));
    InMux I__11612 (
            .O(N__49418),
            .I(N__49278));
    LocalMux I__11611 (
            .O(N__49415),
            .I(N__49267));
    LocalMux I__11610 (
            .O(N__49408),
            .I(N__49267));
    LocalMux I__11609 (
            .O(N__49403),
            .I(N__49267));
    Span4Mux_h I__11608 (
            .O(N__49400),
            .I(N__49267));
    Span4Mux_h I__11607 (
            .O(N__49395),
            .I(N__49267));
    LocalMux I__11606 (
            .O(N__49392),
            .I(N__49264));
    LocalMux I__11605 (
            .O(N__49383),
            .I(N__49257));
    Span4Mux_v I__11604 (
            .O(N__49372),
            .I(N__49257));
    Span4Mux_v I__11603 (
            .O(N__49367),
            .I(N__49257));
    Span4Mux_h I__11602 (
            .O(N__49364),
            .I(N__49250));
    LocalMux I__11601 (
            .O(N__49357),
            .I(N__49250));
    Span4Mux_v I__11600 (
            .O(N__49354),
            .I(N__49250));
    InMux I__11599 (
            .O(N__49353),
            .I(N__49247));
    InMux I__11598 (
            .O(N__49352),
            .I(N__49242));
    InMux I__11597 (
            .O(N__49351),
            .I(N__49242));
    InMux I__11596 (
            .O(N__49350),
            .I(N__49239));
    LocalMux I__11595 (
            .O(N__49343),
            .I(N__49232));
    Span4Mux_h I__11594 (
            .O(N__49340),
            .I(N__49232));
    Span4Mux_h I__11593 (
            .O(N__49337),
            .I(N__49232));
    InMux I__11592 (
            .O(N__49336),
            .I(N__49229));
    InMux I__11591 (
            .O(N__49335),
            .I(N__49224));
    InMux I__11590 (
            .O(N__49334),
            .I(N__49224));
    LocalMux I__11589 (
            .O(N__49329),
            .I(N__49219));
    LocalMux I__11588 (
            .O(N__49322),
            .I(N__49219));
    InMux I__11587 (
            .O(N__49321),
            .I(N__49210));
    InMux I__11586 (
            .O(N__49320),
            .I(N__49210));
    InMux I__11585 (
            .O(N__49319),
            .I(N__49210));
    InMux I__11584 (
            .O(N__49318),
            .I(N__49210));
    LocalMux I__11583 (
            .O(N__49313),
            .I(N__49203));
    Span12Mux_h I__11582 (
            .O(N__49304),
            .I(N__49203));
    LocalMux I__11581 (
            .O(N__49301),
            .I(N__49203));
    Span4Mux_v I__11580 (
            .O(N__49298),
            .I(N__49196));
    LocalMux I__11579 (
            .O(N__49295),
            .I(N__49196));
    LocalMux I__11578 (
            .O(N__49288),
            .I(N__49196));
    LocalMux I__11577 (
            .O(N__49281),
            .I(N__49189));
    LocalMux I__11576 (
            .O(N__49278),
            .I(N__49189));
    Span4Mux_h I__11575 (
            .O(N__49267),
            .I(N__49189));
    Span4Mux_h I__11574 (
            .O(N__49264),
            .I(N__49182));
    Span4Mux_h I__11573 (
            .O(N__49257),
            .I(N__49182));
    Span4Mux_v I__11572 (
            .O(N__49250),
            .I(N__49182));
    LocalMux I__11571 (
            .O(N__49247),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11570 (
            .O(N__49242),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11569 (
            .O(N__49239),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11568 (
            .O(N__49232),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11567 (
            .O(N__49229),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11566 (
            .O(N__49224),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__11565 (
            .O(N__49219),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11564 (
            .O(N__49210),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__11563 (
            .O(N__49203),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11562 (
            .O(N__49196),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11561 (
            .O(N__49189),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11560 (
            .O(N__49182),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__11559 (
            .O(N__49157),
            .I(N__49154));
    LocalMux I__11558 (
            .O(N__49154),
            .I(N__49151));
    Odrv12 I__11557 (
            .O(N__49151),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    ClkMux I__11556 (
            .O(N__49148),
            .I(N__48725));
    ClkMux I__11555 (
            .O(N__49147),
            .I(N__48725));
    ClkMux I__11554 (
            .O(N__49146),
            .I(N__48725));
    ClkMux I__11553 (
            .O(N__49145),
            .I(N__48725));
    ClkMux I__11552 (
            .O(N__49144),
            .I(N__48725));
    ClkMux I__11551 (
            .O(N__49143),
            .I(N__48725));
    ClkMux I__11550 (
            .O(N__49142),
            .I(N__48725));
    ClkMux I__11549 (
            .O(N__49141),
            .I(N__48725));
    ClkMux I__11548 (
            .O(N__49140),
            .I(N__48725));
    ClkMux I__11547 (
            .O(N__49139),
            .I(N__48725));
    ClkMux I__11546 (
            .O(N__49138),
            .I(N__48725));
    ClkMux I__11545 (
            .O(N__49137),
            .I(N__48725));
    ClkMux I__11544 (
            .O(N__49136),
            .I(N__48725));
    ClkMux I__11543 (
            .O(N__49135),
            .I(N__48725));
    ClkMux I__11542 (
            .O(N__49134),
            .I(N__48725));
    ClkMux I__11541 (
            .O(N__49133),
            .I(N__48725));
    ClkMux I__11540 (
            .O(N__49132),
            .I(N__48725));
    ClkMux I__11539 (
            .O(N__49131),
            .I(N__48725));
    ClkMux I__11538 (
            .O(N__49130),
            .I(N__48725));
    ClkMux I__11537 (
            .O(N__49129),
            .I(N__48725));
    ClkMux I__11536 (
            .O(N__49128),
            .I(N__48725));
    ClkMux I__11535 (
            .O(N__49127),
            .I(N__48725));
    ClkMux I__11534 (
            .O(N__49126),
            .I(N__48725));
    ClkMux I__11533 (
            .O(N__49125),
            .I(N__48725));
    ClkMux I__11532 (
            .O(N__49124),
            .I(N__48725));
    ClkMux I__11531 (
            .O(N__49123),
            .I(N__48725));
    ClkMux I__11530 (
            .O(N__49122),
            .I(N__48725));
    ClkMux I__11529 (
            .O(N__49121),
            .I(N__48725));
    ClkMux I__11528 (
            .O(N__49120),
            .I(N__48725));
    ClkMux I__11527 (
            .O(N__49119),
            .I(N__48725));
    ClkMux I__11526 (
            .O(N__49118),
            .I(N__48725));
    ClkMux I__11525 (
            .O(N__49117),
            .I(N__48725));
    ClkMux I__11524 (
            .O(N__49116),
            .I(N__48725));
    ClkMux I__11523 (
            .O(N__49115),
            .I(N__48725));
    ClkMux I__11522 (
            .O(N__49114),
            .I(N__48725));
    ClkMux I__11521 (
            .O(N__49113),
            .I(N__48725));
    ClkMux I__11520 (
            .O(N__49112),
            .I(N__48725));
    ClkMux I__11519 (
            .O(N__49111),
            .I(N__48725));
    ClkMux I__11518 (
            .O(N__49110),
            .I(N__48725));
    ClkMux I__11517 (
            .O(N__49109),
            .I(N__48725));
    ClkMux I__11516 (
            .O(N__49108),
            .I(N__48725));
    ClkMux I__11515 (
            .O(N__49107),
            .I(N__48725));
    ClkMux I__11514 (
            .O(N__49106),
            .I(N__48725));
    ClkMux I__11513 (
            .O(N__49105),
            .I(N__48725));
    ClkMux I__11512 (
            .O(N__49104),
            .I(N__48725));
    ClkMux I__11511 (
            .O(N__49103),
            .I(N__48725));
    ClkMux I__11510 (
            .O(N__49102),
            .I(N__48725));
    ClkMux I__11509 (
            .O(N__49101),
            .I(N__48725));
    ClkMux I__11508 (
            .O(N__49100),
            .I(N__48725));
    ClkMux I__11507 (
            .O(N__49099),
            .I(N__48725));
    ClkMux I__11506 (
            .O(N__49098),
            .I(N__48725));
    ClkMux I__11505 (
            .O(N__49097),
            .I(N__48725));
    ClkMux I__11504 (
            .O(N__49096),
            .I(N__48725));
    ClkMux I__11503 (
            .O(N__49095),
            .I(N__48725));
    ClkMux I__11502 (
            .O(N__49094),
            .I(N__48725));
    ClkMux I__11501 (
            .O(N__49093),
            .I(N__48725));
    ClkMux I__11500 (
            .O(N__49092),
            .I(N__48725));
    ClkMux I__11499 (
            .O(N__49091),
            .I(N__48725));
    ClkMux I__11498 (
            .O(N__49090),
            .I(N__48725));
    ClkMux I__11497 (
            .O(N__49089),
            .I(N__48725));
    ClkMux I__11496 (
            .O(N__49088),
            .I(N__48725));
    ClkMux I__11495 (
            .O(N__49087),
            .I(N__48725));
    ClkMux I__11494 (
            .O(N__49086),
            .I(N__48725));
    ClkMux I__11493 (
            .O(N__49085),
            .I(N__48725));
    ClkMux I__11492 (
            .O(N__49084),
            .I(N__48725));
    ClkMux I__11491 (
            .O(N__49083),
            .I(N__48725));
    ClkMux I__11490 (
            .O(N__49082),
            .I(N__48725));
    ClkMux I__11489 (
            .O(N__49081),
            .I(N__48725));
    ClkMux I__11488 (
            .O(N__49080),
            .I(N__48725));
    ClkMux I__11487 (
            .O(N__49079),
            .I(N__48725));
    ClkMux I__11486 (
            .O(N__49078),
            .I(N__48725));
    ClkMux I__11485 (
            .O(N__49077),
            .I(N__48725));
    ClkMux I__11484 (
            .O(N__49076),
            .I(N__48725));
    ClkMux I__11483 (
            .O(N__49075),
            .I(N__48725));
    ClkMux I__11482 (
            .O(N__49074),
            .I(N__48725));
    ClkMux I__11481 (
            .O(N__49073),
            .I(N__48725));
    ClkMux I__11480 (
            .O(N__49072),
            .I(N__48725));
    ClkMux I__11479 (
            .O(N__49071),
            .I(N__48725));
    ClkMux I__11478 (
            .O(N__49070),
            .I(N__48725));
    ClkMux I__11477 (
            .O(N__49069),
            .I(N__48725));
    ClkMux I__11476 (
            .O(N__49068),
            .I(N__48725));
    ClkMux I__11475 (
            .O(N__49067),
            .I(N__48725));
    ClkMux I__11474 (
            .O(N__49066),
            .I(N__48725));
    ClkMux I__11473 (
            .O(N__49065),
            .I(N__48725));
    ClkMux I__11472 (
            .O(N__49064),
            .I(N__48725));
    ClkMux I__11471 (
            .O(N__49063),
            .I(N__48725));
    ClkMux I__11470 (
            .O(N__49062),
            .I(N__48725));
    ClkMux I__11469 (
            .O(N__49061),
            .I(N__48725));
    ClkMux I__11468 (
            .O(N__49060),
            .I(N__48725));
    ClkMux I__11467 (
            .O(N__49059),
            .I(N__48725));
    ClkMux I__11466 (
            .O(N__49058),
            .I(N__48725));
    ClkMux I__11465 (
            .O(N__49057),
            .I(N__48725));
    ClkMux I__11464 (
            .O(N__49056),
            .I(N__48725));
    ClkMux I__11463 (
            .O(N__49055),
            .I(N__48725));
    ClkMux I__11462 (
            .O(N__49054),
            .I(N__48725));
    ClkMux I__11461 (
            .O(N__49053),
            .I(N__48725));
    ClkMux I__11460 (
            .O(N__49052),
            .I(N__48725));
    ClkMux I__11459 (
            .O(N__49051),
            .I(N__48725));
    ClkMux I__11458 (
            .O(N__49050),
            .I(N__48725));
    ClkMux I__11457 (
            .O(N__49049),
            .I(N__48725));
    ClkMux I__11456 (
            .O(N__49048),
            .I(N__48725));
    ClkMux I__11455 (
            .O(N__49047),
            .I(N__48725));
    ClkMux I__11454 (
            .O(N__49046),
            .I(N__48725));
    ClkMux I__11453 (
            .O(N__49045),
            .I(N__48725));
    ClkMux I__11452 (
            .O(N__49044),
            .I(N__48725));
    ClkMux I__11451 (
            .O(N__49043),
            .I(N__48725));
    ClkMux I__11450 (
            .O(N__49042),
            .I(N__48725));
    ClkMux I__11449 (
            .O(N__49041),
            .I(N__48725));
    ClkMux I__11448 (
            .O(N__49040),
            .I(N__48725));
    ClkMux I__11447 (
            .O(N__49039),
            .I(N__48725));
    ClkMux I__11446 (
            .O(N__49038),
            .I(N__48725));
    ClkMux I__11445 (
            .O(N__49037),
            .I(N__48725));
    ClkMux I__11444 (
            .O(N__49036),
            .I(N__48725));
    ClkMux I__11443 (
            .O(N__49035),
            .I(N__48725));
    ClkMux I__11442 (
            .O(N__49034),
            .I(N__48725));
    ClkMux I__11441 (
            .O(N__49033),
            .I(N__48725));
    ClkMux I__11440 (
            .O(N__49032),
            .I(N__48725));
    ClkMux I__11439 (
            .O(N__49031),
            .I(N__48725));
    ClkMux I__11438 (
            .O(N__49030),
            .I(N__48725));
    ClkMux I__11437 (
            .O(N__49029),
            .I(N__48725));
    ClkMux I__11436 (
            .O(N__49028),
            .I(N__48725));
    ClkMux I__11435 (
            .O(N__49027),
            .I(N__48725));
    ClkMux I__11434 (
            .O(N__49026),
            .I(N__48725));
    ClkMux I__11433 (
            .O(N__49025),
            .I(N__48725));
    ClkMux I__11432 (
            .O(N__49024),
            .I(N__48725));
    ClkMux I__11431 (
            .O(N__49023),
            .I(N__48725));
    ClkMux I__11430 (
            .O(N__49022),
            .I(N__48725));
    ClkMux I__11429 (
            .O(N__49021),
            .I(N__48725));
    ClkMux I__11428 (
            .O(N__49020),
            .I(N__48725));
    ClkMux I__11427 (
            .O(N__49019),
            .I(N__48725));
    ClkMux I__11426 (
            .O(N__49018),
            .I(N__48725));
    ClkMux I__11425 (
            .O(N__49017),
            .I(N__48725));
    ClkMux I__11424 (
            .O(N__49016),
            .I(N__48725));
    ClkMux I__11423 (
            .O(N__49015),
            .I(N__48725));
    ClkMux I__11422 (
            .O(N__49014),
            .I(N__48725));
    ClkMux I__11421 (
            .O(N__49013),
            .I(N__48725));
    ClkMux I__11420 (
            .O(N__49012),
            .I(N__48725));
    ClkMux I__11419 (
            .O(N__49011),
            .I(N__48725));
    ClkMux I__11418 (
            .O(N__49010),
            .I(N__48725));
    ClkMux I__11417 (
            .O(N__49009),
            .I(N__48725));
    ClkMux I__11416 (
            .O(N__49008),
            .I(N__48725));
    GlobalMux I__11415 (
            .O(N__48725),
            .I(clk_100mhz_0));
    CEMux I__11414 (
            .O(N__48722),
            .I(N__48689));
    CEMux I__11413 (
            .O(N__48721),
            .I(N__48689));
    CEMux I__11412 (
            .O(N__48720),
            .I(N__48689));
    CEMux I__11411 (
            .O(N__48719),
            .I(N__48689));
    CEMux I__11410 (
            .O(N__48718),
            .I(N__48689));
    CEMux I__11409 (
            .O(N__48717),
            .I(N__48689));
    CEMux I__11408 (
            .O(N__48716),
            .I(N__48689));
    CEMux I__11407 (
            .O(N__48715),
            .I(N__48689));
    CEMux I__11406 (
            .O(N__48714),
            .I(N__48689));
    CEMux I__11405 (
            .O(N__48713),
            .I(N__48689));
    CEMux I__11404 (
            .O(N__48712),
            .I(N__48689));
    GlobalMux I__11403 (
            .O(N__48689),
            .I(N__48686));
    gio2CtrlBuf I__11402 (
            .O(N__48686),
            .I(\phase_controller_inst2.stoper_hc.un1_start_g ));
    InMux I__11401 (
            .O(N__48683),
            .I(N__48677));
    InMux I__11400 (
            .O(N__48682),
            .I(N__48674));
    InMux I__11399 (
            .O(N__48681),
            .I(N__48671));
    InMux I__11398 (
            .O(N__48680),
            .I(N__48668));
    LocalMux I__11397 (
            .O(N__48677),
            .I(N__48665));
    LocalMux I__11396 (
            .O(N__48674),
            .I(N__48662));
    LocalMux I__11395 (
            .O(N__48671),
            .I(N__48659));
    LocalMux I__11394 (
            .O(N__48668),
            .I(N__48560));
    Glb2LocalMux I__11393 (
            .O(N__48665),
            .I(N__48227));
    Glb2LocalMux I__11392 (
            .O(N__48662),
            .I(N__48227));
    Glb2LocalMux I__11391 (
            .O(N__48659),
            .I(N__48227));
    SRMux I__11390 (
            .O(N__48658),
            .I(N__48227));
    SRMux I__11389 (
            .O(N__48657),
            .I(N__48227));
    SRMux I__11388 (
            .O(N__48656),
            .I(N__48227));
    SRMux I__11387 (
            .O(N__48655),
            .I(N__48227));
    SRMux I__11386 (
            .O(N__48654),
            .I(N__48227));
    SRMux I__11385 (
            .O(N__48653),
            .I(N__48227));
    SRMux I__11384 (
            .O(N__48652),
            .I(N__48227));
    SRMux I__11383 (
            .O(N__48651),
            .I(N__48227));
    SRMux I__11382 (
            .O(N__48650),
            .I(N__48227));
    SRMux I__11381 (
            .O(N__48649),
            .I(N__48227));
    SRMux I__11380 (
            .O(N__48648),
            .I(N__48227));
    SRMux I__11379 (
            .O(N__48647),
            .I(N__48227));
    SRMux I__11378 (
            .O(N__48646),
            .I(N__48227));
    SRMux I__11377 (
            .O(N__48645),
            .I(N__48227));
    SRMux I__11376 (
            .O(N__48644),
            .I(N__48227));
    SRMux I__11375 (
            .O(N__48643),
            .I(N__48227));
    SRMux I__11374 (
            .O(N__48642),
            .I(N__48227));
    SRMux I__11373 (
            .O(N__48641),
            .I(N__48227));
    SRMux I__11372 (
            .O(N__48640),
            .I(N__48227));
    SRMux I__11371 (
            .O(N__48639),
            .I(N__48227));
    SRMux I__11370 (
            .O(N__48638),
            .I(N__48227));
    SRMux I__11369 (
            .O(N__48637),
            .I(N__48227));
    SRMux I__11368 (
            .O(N__48636),
            .I(N__48227));
    SRMux I__11367 (
            .O(N__48635),
            .I(N__48227));
    SRMux I__11366 (
            .O(N__48634),
            .I(N__48227));
    SRMux I__11365 (
            .O(N__48633),
            .I(N__48227));
    SRMux I__11364 (
            .O(N__48632),
            .I(N__48227));
    SRMux I__11363 (
            .O(N__48631),
            .I(N__48227));
    SRMux I__11362 (
            .O(N__48630),
            .I(N__48227));
    SRMux I__11361 (
            .O(N__48629),
            .I(N__48227));
    SRMux I__11360 (
            .O(N__48628),
            .I(N__48227));
    SRMux I__11359 (
            .O(N__48627),
            .I(N__48227));
    SRMux I__11358 (
            .O(N__48626),
            .I(N__48227));
    SRMux I__11357 (
            .O(N__48625),
            .I(N__48227));
    SRMux I__11356 (
            .O(N__48624),
            .I(N__48227));
    SRMux I__11355 (
            .O(N__48623),
            .I(N__48227));
    SRMux I__11354 (
            .O(N__48622),
            .I(N__48227));
    SRMux I__11353 (
            .O(N__48621),
            .I(N__48227));
    SRMux I__11352 (
            .O(N__48620),
            .I(N__48227));
    SRMux I__11351 (
            .O(N__48619),
            .I(N__48227));
    SRMux I__11350 (
            .O(N__48618),
            .I(N__48227));
    SRMux I__11349 (
            .O(N__48617),
            .I(N__48227));
    SRMux I__11348 (
            .O(N__48616),
            .I(N__48227));
    SRMux I__11347 (
            .O(N__48615),
            .I(N__48227));
    SRMux I__11346 (
            .O(N__48614),
            .I(N__48227));
    SRMux I__11345 (
            .O(N__48613),
            .I(N__48227));
    SRMux I__11344 (
            .O(N__48612),
            .I(N__48227));
    SRMux I__11343 (
            .O(N__48611),
            .I(N__48227));
    SRMux I__11342 (
            .O(N__48610),
            .I(N__48227));
    SRMux I__11341 (
            .O(N__48609),
            .I(N__48227));
    SRMux I__11340 (
            .O(N__48608),
            .I(N__48227));
    SRMux I__11339 (
            .O(N__48607),
            .I(N__48227));
    SRMux I__11338 (
            .O(N__48606),
            .I(N__48227));
    SRMux I__11337 (
            .O(N__48605),
            .I(N__48227));
    SRMux I__11336 (
            .O(N__48604),
            .I(N__48227));
    SRMux I__11335 (
            .O(N__48603),
            .I(N__48227));
    SRMux I__11334 (
            .O(N__48602),
            .I(N__48227));
    SRMux I__11333 (
            .O(N__48601),
            .I(N__48227));
    SRMux I__11332 (
            .O(N__48600),
            .I(N__48227));
    SRMux I__11331 (
            .O(N__48599),
            .I(N__48227));
    SRMux I__11330 (
            .O(N__48598),
            .I(N__48227));
    SRMux I__11329 (
            .O(N__48597),
            .I(N__48227));
    SRMux I__11328 (
            .O(N__48596),
            .I(N__48227));
    SRMux I__11327 (
            .O(N__48595),
            .I(N__48227));
    SRMux I__11326 (
            .O(N__48594),
            .I(N__48227));
    SRMux I__11325 (
            .O(N__48593),
            .I(N__48227));
    SRMux I__11324 (
            .O(N__48592),
            .I(N__48227));
    SRMux I__11323 (
            .O(N__48591),
            .I(N__48227));
    SRMux I__11322 (
            .O(N__48590),
            .I(N__48227));
    SRMux I__11321 (
            .O(N__48589),
            .I(N__48227));
    SRMux I__11320 (
            .O(N__48588),
            .I(N__48227));
    SRMux I__11319 (
            .O(N__48587),
            .I(N__48227));
    SRMux I__11318 (
            .O(N__48586),
            .I(N__48227));
    SRMux I__11317 (
            .O(N__48585),
            .I(N__48227));
    SRMux I__11316 (
            .O(N__48584),
            .I(N__48227));
    SRMux I__11315 (
            .O(N__48583),
            .I(N__48227));
    SRMux I__11314 (
            .O(N__48582),
            .I(N__48227));
    SRMux I__11313 (
            .O(N__48581),
            .I(N__48227));
    SRMux I__11312 (
            .O(N__48580),
            .I(N__48227));
    SRMux I__11311 (
            .O(N__48579),
            .I(N__48227));
    SRMux I__11310 (
            .O(N__48578),
            .I(N__48227));
    SRMux I__11309 (
            .O(N__48577),
            .I(N__48227));
    SRMux I__11308 (
            .O(N__48576),
            .I(N__48227));
    SRMux I__11307 (
            .O(N__48575),
            .I(N__48227));
    SRMux I__11306 (
            .O(N__48574),
            .I(N__48227));
    SRMux I__11305 (
            .O(N__48573),
            .I(N__48227));
    SRMux I__11304 (
            .O(N__48572),
            .I(N__48227));
    SRMux I__11303 (
            .O(N__48571),
            .I(N__48227));
    SRMux I__11302 (
            .O(N__48570),
            .I(N__48227));
    SRMux I__11301 (
            .O(N__48569),
            .I(N__48227));
    SRMux I__11300 (
            .O(N__48568),
            .I(N__48227));
    SRMux I__11299 (
            .O(N__48567),
            .I(N__48227));
    SRMux I__11298 (
            .O(N__48566),
            .I(N__48227));
    SRMux I__11297 (
            .O(N__48565),
            .I(N__48227));
    SRMux I__11296 (
            .O(N__48564),
            .I(N__48227));
    SRMux I__11295 (
            .O(N__48563),
            .I(N__48227));
    Glb2LocalMux I__11294 (
            .O(N__48560),
            .I(N__48227));
    SRMux I__11293 (
            .O(N__48559),
            .I(N__48227));
    SRMux I__11292 (
            .O(N__48558),
            .I(N__48227));
    SRMux I__11291 (
            .O(N__48557),
            .I(N__48227));
    SRMux I__11290 (
            .O(N__48556),
            .I(N__48227));
    SRMux I__11289 (
            .O(N__48555),
            .I(N__48227));
    SRMux I__11288 (
            .O(N__48554),
            .I(N__48227));
    SRMux I__11287 (
            .O(N__48553),
            .I(N__48227));
    SRMux I__11286 (
            .O(N__48552),
            .I(N__48227));
    SRMux I__11285 (
            .O(N__48551),
            .I(N__48227));
    SRMux I__11284 (
            .O(N__48550),
            .I(N__48227));
    SRMux I__11283 (
            .O(N__48549),
            .I(N__48227));
    SRMux I__11282 (
            .O(N__48548),
            .I(N__48227));
    SRMux I__11281 (
            .O(N__48547),
            .I(N__48227));
    SRMux I__11280 (
            .O(N__48546),
            .I(N__48227));
    SRMux I__11279 (
            .O(N__48545),
            .I(N__48227));
    SRMux I__11278 (
            .O(N__48544),
            .I(N__48227));
    SRMux I__11277 (
            .O(N__48543),
            .I(N__48227));
    SRMux I__11276 (
            .O(N__48542),
            .I(N__48227));
    SRMux I__11275 (
            .O(N__48541),
            .I(N__48227));
    SRMux I__11274 (
            .O(N__48540),
            .I(N__48227));
    SRMux I__11273 (
            .O(N__48539),
            .I(N__48227));
    SRMux I__11272 (
            .O(N__48538),
            .I(N__48227));
    SRMux I__11271 (
            .O(N__48537),
            .I(N__48227));
    SRMux I__11270 (
            .O(N__48536),
            .I(N__48227));
    SRMux I__11269 (
            .O(N__48535),
            .I(N__48227));
    SRMux I__11268 (
            .O(N__48534),
            .I(N__48227));
    SRMux I__11267 (
            .O(N__48533),
            .I(N__48227));
    SRMux I__11266 (
            .O(N__48532),
            .I(N__48227));
    SRMux I__11265 (
            .O(N__48531),
            .I(N__48227));
    SRMux I__11264 (
            .O(N__48530),
            .I(N__48227));
    SRMux I__11263 (
            .O(N__48529),
            .I(N__48227));
    SRMux I__11262 (
            .O(N__48528),
            .I(N__48227));
    SRMux I__11261 (
            .O(N__48527),
            .I(N__48227));
    SRMux I__11260 (
            .O(N__48526),
            .I(N__48227));
    SRMux I__11259 (
            .O(N__48525),
            .I(N__48227));
    SRMux I__11258 (
            .O(N__48524),
            .I(N__48227));
    SRMux I__11257 (
            .O(N__48523),
            .I(N__48227));
    SRMux I__11256 (
            .O(N__48522),
            .I(N__48227));
    SRMux I__11255 (
            .O(N__48521),
            .I(N__48227));
    SRMux I__11254 (
            .O(N__48520),
            .I(N__48227));
    SRMux I__11253 (
            .O(N__48519),
            .I(N__48227));
    SRMux I__11252 (
            .O(N__48518),
            .I(N__48227));
    SRMux I__11251 (
            .O(N__48517),
            .I(N__48227));
    SRMux I__11250 (
            .O(N__48516),
            .I(N__48227));
    GlobalMux I__11249 (
            .O(N__48227),
            .I(N__48224));
    gio2CtrlBuf I__11248 (
            .O(N__48224),
            .I(red_c_g));
    InMux I__11247 (
            .O(N__48221),
            .I(N__48218));
    LocalMux I__11246 (
            .O(N__48218),
            .I(N__48215));
    Span4Mux_v I__11245 (
            .O(N__48215),
            .I(N__48211));
    InMux I__11244 (
            .O(N__48214),
            .I(N__48208));
    Odrv4 I__11243 (
            .O(N__48211),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__11242 (
            .O(N__48208),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    CascadeMux I__11241 (
            .O(N__48203),
            .I(elapsed_time_ns_1_RNI57CN9_0_18_cascade_));
    InMux I__11240 (
            .O(N__48200),
            .I(N__48194));
    InMux I__11239 (
            .O(N__48199),
            .I(N__48194));
    LocalMux I__11238 (
            .O(N__48194),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    InMux I__11237 (
            .O(N__48191),
            .I(N__48188));
    LocalMux I__11236 (
            .O(N__48188),
            .I(N__48185));
    Span4Mux_v I__11235 (
            .O(N__48185),
            .I(N__48182));
    Odrv4 I__11234 (
            .O(N__48182),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt26 ));
    InMux I__11233 (
            .O(N__48179),
            .I(N__48173));
    InMux I__11232 (
            .O(N__48178),
            .I(N__48173));
    LocalMux I__11231 (
            .O(N__48173),
            .I(N__48169));
    InMux I__11230 (
            .O(N__48172),
            .I(N__48165));
    Span4Mux_v I__11229 (
            .O(N__48169),
            .I(N__48162));
    InMux I__11228 (
            .O(N__48168),
            .I(N__48159));
    LocalMux I__11227 (
            .O(N__48165),
            .I(N__48152));
    Span4Mux_v I__11226 (
            .O(N__48162),
            .I(N__48152));
    LocalMux I__11225 (
            .O(N__48159),
            .I(N__48152));
    Odrv4 I__11224 (
            .O(N__48152),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__11223 (
            .O(N__48149),
            .I(N__48144));
    InMux I__11222 (
            .O(N__48148),
            .I(N__48140));
    InMux I__11221 (
            .O(N__48147),
            .I(N__48137));
    LocalMux I__11220 (
            .O(N__48144),
            .I(N__48134));
    InMux I__11219 (
            .O(N__48143),
            .I(N__48131));
    LocalMux I__11218 (
            .O(N__48140),
            .I(N__48126));
    LocalMux I__11217 (
            .O(N__48137),
            .I(N__48126));
    Span4Mux_h I__11216 (
            .O(N__48134),
            .I(N__48121));
    LocalMux I__11215 (
            .O(N__48131),
            .I(N__48121));
    Span4Mux_v I__11214 (
            .O(N__48126),
            .I(N__48118));
    Odrv4 I__11213 (
            .O(N__48121),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__11212 (
            .O(N__48118),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    CascadeMux I__11211 (
            .O(N__48113),
            .I(N__48108));
    InMux I__11210 (
            .O(N__48112),
            .I(N__48104));
    InMux I__11209 (
            .O(N__48111),
            .I(N__48101));
    InMux I__11208 (
            .O(N__48108),
            .I(N__48098));
    InMux I__11207 (
            .O(N__48107),
            .I(N__48095));
    LocalMux I__11206 (
            .O(N__48104),
            .I(N__48092));
    LocalMux I__11205 (
            .O(N__48101),
            .I(N__48087));
    LocalMux I__11204 (
            .O(N__48098),
            .I(N__48087));
    LocalMux I__11203 (
            .O(N__48095),
            .I(N__48084));
    Span4Mux_v I__11202 (
            .O(N__48092),
            .I(N__48079));
    Span4Mux_v I__11201 (
            .O(N__48087),
            .I(N__48079));
    Odrv12 I__11200 (
            .O(N__48084),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv4 I__11199 (
            .O(N__48079),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__11198 (
            .O(N__48074),
            .I(N__48067));
    InMux I__11197 (
            .O(N__48073),
            .I(N__48067));
    InMux I__11196 (
            .O(N__48072),
            .I(N__48063));
    LocalMux I__11195 (
            .O(N__48067),
            .I(N__48060));
    InMux I__11194 (
            .O(N__48066),
            .I(N__48057));
    LocalMux I__11193 (
            .O(N__48063),
            .I(N__48054));
    Span4Mux_v I__11192 (
            .O(N__48060),
            .I(N__48049));
    LocalMux I__11191 (
            .O(N__48057),
            .I(N__48049));
    Odrv4 I__11190 (
            .O(N__48054),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv4 I__11189 (
            .O(N__48049),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__11188 (
            .O(N__48044),
            .I(N__48041));
    LocalMux I__11187 (
            .O(N__48041),
            .I(N__48038));
    Odrv4 I__11186 (
            .O(N__48038),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ));
    InMux I__11185 (
            .O(N__48035),
            .I(N__48032));
    LocalMux I__11184 (
            .O(N__48032),
            .I(N__48029));
    Odrv4 I__11183 (
            .O(N__48029),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    CascadeMux I__11182 (
            .O(N__48026),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_ ));
    CascadeMux I__11181 (
            .O(N__48023),
            .I(N__48020));
    InMux I__11180 (
            .O(N__48020),
            .I(N__48017));
    LocalMux I__11179 (
            .O(N__48017),
            .I(N__48014));
    Span4Mux_h I__11178 (
            .O(N__48014),
            .I(N__48011));
    Span4Mux_h I__11177 (
            .O(N__48011),
            .I(N__48008));
    Odrv4 I__11176 (
            .O(N__48008),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    InMux I__11175 (
            .O(N__48005),
            .I(N__48000));
    InMux I__11174 (
            .O(N__48004),
            .I(N__47995));
    InMux I__11173 (
            .O(N__48003),
            .I(N__47995));
    LocalMux I__11172 (
            .O(N__48000),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__11171 (
            .O(N__47995),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__11170 (
            .O(N__47990),
            .I(N__47985));
    InMux I__11169 (
            .O(N__47989),
            .I(N__47980));
    InMux I__11168 (
            .O(N__47988),
            .I(N__47980));
    LocalMux I__11167 (
            .O(N__47985),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__11166 (
            .O(N__47980),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    CascadeMux I__11165 (
            .O(N__47975),
            .I(N__47972));
    InMux I__11164 (
            .O(N__47972),
            .I(N__47969));
    LocalMux I__11163 (
            .O(N__47969),
            .I(N__47966));
    Span4Mux_v I__11162 (
            .O(N__47966),
            .I(N__47963));
    Odrv4 I__11161 (
            .O(N__47963),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ));
    InMux I__11160 (
            .O(N__47960),
            .I(N__47955));
    InMux I__11159 (
            .O(N__47959),
            .I(N__47952));
    InMux I__11158 (
            .O(N__47958),
            .I(N__47949));
    LocalMux I__11157 (
            .O(N__47955),
            .I(N__47945));
    LocalMux I__11156 (
            .O(N__47952),
            .I(N__47942));
    LocalMux I__11155 (
            .O(N__47949),
            .I(N__47939));
    CascadeMux I__11154 (
            .O(N__47948),
            .I(N__47936));
    Span4Mux_h I__11153 (
            .O(N__47945),
            .I(N__47931));
    Span4Mux_h I__11152 (
            .O(N__47942),
            .I(N__47931));
    Span4Mux_h I__11151 (
            .O(N__47939),
            .I(N__47928));
    InMux I__11150 (
            .O(N__47936),
            .I(N__47925));
    Odrv4 I__11149 (
            .O(N__47931),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__11148 (
            .O(N__47928),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    LocalMux I__11147 (
            .O(N__47925),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__11146 (
            .O(N__47918),
            .I(N__47915));
    LocalMux I__11145 (
            .O(N__47915),
            .I(N__47910));
    InMux I__11144 (
            .O(N__47914),
            .I(N__47907));
    InMux I__11143 (
            .O(N__47913),
            .I(N__47904));
    Span4Mux_h I__11142 (
            .O(N__47910),
            .I(N__47901));
    LocalMux I__11141 (
            .O(N__47907),
            .I(N__47898));
    LocalMux I__11140 (
            .O(N__47904),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv4 I__11139 (
            .O(N__47901),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv4 I__11138 (
            .O(N__47898),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    InMux I__11137 (
            .O(N__47891),
            .I(N__47887));
    InMux I__11136 (
            .O(N__47890),
            .I(N__47882));
    LocalMux I__11135 (
            .O(N__47887),
            .I(N__47879));
    InMux I__11134 (
            .O(N__47886),
            .I(N__47876));
    InMux I__11133 (
            .O(N__47885),
            .I(N__47873));
    LocalMux I__11132 (
            .O(N__47882),
            .I(N__47870));
    Span4Mux_h I__11131 (
            .O(N__47879),
            .I(N__47867));
    LocalMux I__11130 (
            .O(N__47876),
            .I(N__47864));
    LocalMux I__11129 (
            .O(N__47873),
            .I(N__47861));
    Odrv12 I__11128 (
            .O(N__47870),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__11127 (
            .O(N__47867),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__11126 (
            .O(N__47864),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__11125 (
            .O(N__47861),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__11124 (
            .O(N__47852),
            .I(N__47845));
    InMux I__11123 (
            .O(N__47851),
            .I(N__47845));
    InMux I__11122 (
            .O(N__47850),
            .I(N__47841));
    LocalMux I__11121 (
            .O(N__47845),
            .I(N__47838));
    InMux I__11120 (
            .O(N__47844),
            .I(N__47835));
    LocalMux I__11119 (
            .O(N__47841),
            .I(N__47832));
    Span4Mux_h I__11118 (
            .O(N__47838),
            .I(N__47829));
    LocalMux I__11117 (
            .O(N__47835),
            .I(N__47826));
    Span4Mux_h I__11116 (
            .O(N__47832),
            .I(N__47823));
    Span4Mux_v I__11115 (
            .O(N__47829),
            .I(N__47820));
    Span4Mux_h I__11114 (
            .O(N__47826),
            .I(N__47817));
    Odrv4 I__11113 (
            .O(N__47823),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__11112 (
            .O(N__47820),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__11111 (
            .O(N__47817),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__11110 (
            .O(N__47810),
            .I(N__47805));
    InMux I__11109 (
            .O(N__47809),
            .I(N__47802));
    InMux I__11108 (
            .O(N__47808),
            .I(N__47798));
    LocalMux I__11107 (
            .O(N__47805),
            .I(N__47793));
    LocalMux I__11106 (
            .O(N__47802),
            .I(N__47793));
    InMux I__11105 (
            .O(N__47801),
            .I(N__47790));
    LocalMux I__11104 (
            .O(N__47798),
            .I(N__47787));
    Span4Mux_v I__11103 (
            .O(N__47793),
            .I(N__47784));
    LocalMux I__11102 (
            .O(N__47790),
            .I(N__47781));
    Odrv4 I__11101 (
            .O(N__47787),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__11100 (
            .O(N__47784),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__11099 (
            .O(N__47781),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__11098 (
            .O(N__47774),
            .I(N__47771));
    LocalMux I__11097 (
            .O(N__47771),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    InMux I__11096 (
            .O(N__47768),
            .I(N__47765));
    LocalMux I__11095 (
            .O(N__47765),
            .I(N__47761));
    InMux I__11094 (
            .O(N__47764),
            .I(N__47758));
    Span4Mux_h I__11093 (
            .O(N__47761),
            .I(N__47753));
    LocalMux I__11092 (
            .O(N__47758),
            .I(N__47750));
    InMux I__11091 (
            .O(N__47757),
            .I(N__47745));
    InMux I__11090 (
            .O(N__47756),
            .I(N__47745));
    Odrv4 I__11089 (
            .O(N__47753),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    Odrv4 I__11088 (
            .O(N__47750),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__11087 (
            .O(N__47745),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__11086 (
            .O(N__47738),
            .I(N__47735));
    LocalMux I__11085 (
            .O(N__47735),
            .I(N__47732));
    Span4Mux_h I__11084 (
            .O(N__47732),
            .I(N__47729));
    Odrv4 I__11083 (
            .O(N__47729),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__11082 (
            .O(N__47726),
            .I(N__47723));
    InMux I__11081 (
            .O(N__47723),
            .I(N__47717));
    InMux I__11080 (
            .O(N__47722),
            .I(N__47717));
    LocalMux I__11079 (
            .O(N__47717),
            .I(N__47714));
    Odrv4 I__11078 (
            .O(N__47714),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    InMux I__11077 (
            .O(N__47711),
            .I(N__47708));
    LocalMux I__11076 (
            .O(N__47708),
            .I(N__47704));
    InMux I__11075 (
            .O(N__47707),
            .I(N__47700));
    Span12Mux_v I__11074 (
            .O(N__47704),
            .I(N__47697));
    InMux I__11073 (
            .O(N__47703),
            .I(N__47694));
    LocalMux I__11072 (
            .O(N__47700),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv12 I__11071 (
            .O(N__47697),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    LocalMux I__11070 (
            .O(N__47694),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    InMux I__11069 (
            .O(N__47687),
            .I(N__47683));
    InMux I__11068 (
            .O(N__47686),
            .I(N__47680));
    LocalMux I__11067 (
            .O(N__47683),
            .I(N__47675));
    LocalMux I__11066 (
            .O(N__47680),
            .I(N__47672));
    InMux I__11065 (
            .O(N__47679),
            .I(N__47669));
    CascadeMux I__11064 (
            .O(N__47678),
            .I(N__47666));
    Span4Mux_h I__11063 (
            .O(N__47675),
            .I(N__47663));
    Span4Mux_v I__11062 (
            .O(N__47672),
            .I(N__47658));
    LocalMux I__11061 (
            .O(N__47669),
            .I(N__47658));
    InMux I__11060 (
            .O(N__47666),
            .I(N__47655));
    Odrv4 I__11059 (
            .O(N__47663),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv4 I__11058 (
            .O(N__47658),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    LocalMux I__11057 (
            .O(N__47655),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__11056 (
            .O(N__47648),
            .I(N__47642));
    InMux I__11055 (
            .O(N__47647),
            .I(N__47642));
    LocalMux I__11054 (
            .O(N__47642),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    InMux I__11053 (
            .O(N__47639),
            .I(N__47636));
    LocalMux I__11052 (
            .O(N__47636),
            .I(N__47632));
    InMux I__11051 (
            .O(N__47635),
            .I(N__47628));
    Span4Mux_v I__11050 (
            .O(N__47632),
            .I(N__47625));
    InMux I__11049 (
            .O(N__47631),
            .I(N__47622));
    LocalMux I__11048 (
            .O(N__47628),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    Odrv4 I__11047 (
            .O(N__47625),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    LocalMux I__11046 (
            .O(N__47622),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    CascadeMux I__11045 (
            .O(N__47615),
            .I(N__47612));
    InMux I__11044 (
            .O(N__47612),
            .I(N__47609));
    LocalMux I__11043 (
            .O(N__47609),
            .I(N__47606));
    Odrv4 I__11042 (
            .O(N__47606),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__11041 (
            .O(N__47603),
            .I(N__47600));
    LocalMux I__11040 (
            .O(N__47600),
            .I(N__47596));
    InMux I__11039 (
            .O(N__47599),
            .I(N__47592));
    Span12Mux_h I__11038 (
            .O(N__47596),
            .I(N__47589));
    InMux I__11037 (
            .O(N__47595),
            .I(N__47586));
    LocalMux I__11036 (
            .O(N__47592),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    Odrv12 I__11035 (
            .O(N__47589),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__11034 (
            .O(N__47586),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    InMux I__11033 (
            .O(N__47579),
            .I(N__47573));
    InMux I__11032 (
            .O(N__47578),
            .I(N__47573));
    LocalMux I__11031 (
            .O(N__47573),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    InMux I__11030 (
            .O(N__47570),
            .I(N__47564));
    InMux I__11029 (
            .O(N__47569),
            .I(N__47564));
    LocalMux I__11028 (
            .O(N__47564),
            .I(N__47561));
    Odrv12 I__11027 (
            .O(N__47561),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__11026 (
            .O(N__47558),
            .I(N__47555));
    InMux I__11025 (
            .O(N__47555),
            .I(N__47552));
    LocalMux I__11024 (
            .O(N__47552),
            .I(N__47549));
    Span4Mux_h I__11023 (
            .O(N__47549),
            .I(N__47546));
    Odrv4 I__11022 (
            .O(N__47546),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    InMux I__11021 (
            .O(N__47543),
            .I(N__47538));
    InMux I__11020 (
            .O(N__47542),
            .I(N__47533));
    InMux I__11019 (
            .O(N__47541),
            .I(N__47533));
    LocalMux I__11018 (
            .O(N__47538),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__11017 (
            .O(N__47533),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__11016 (
            .O(N__47528),
            .I(N__47524));
    InMux I__11015 (
            .O(N__47527),
            .I(N__47520));
    InMux I__11014 (
            .O(N__47524),
            .I(N__47515));
    InMux I__11013 (
            .O(N__47523),
            .I(N__47515));
    LocalMux I__11012 (
            .O(N__47520),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__11011 (
            .O(N__47515),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__11010 (
            .O(N__47510),
            .I(N__47507));
    LocalMux I__11009 (
            .O(N__47507),
            .I(N__47504));
    Odrv4 I__11008 (
            .O(N__47504),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    InMux I__11007 (
            .O(N__47501),
            .I(N__47497));
    InMux I__11006 (
            .O(N__47500),
            .I(N__47494));
    LocalMux I__11005 (
            .O(N__47497),
            .I(N__47490));
    LocalMux I__11004 (
            .O(N__47494),
            .I(N__47487));
    InMux I__11003 (
            .O(N__47493),
            .I(N__47484));
    Span4Mux_h I__11002 (
            .O(N__47490),
            .I(N__47479));
    Span4Mux_h I__11001 (
            .O(N__47487),
            .I(N__47479));
    LocalMux I__11000 (
            .O(N__47484),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    Odrv4 I__10999 (
            .O(N__47479),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    CascadeMux I__10998 (
            .O(N__47474),
            .I(N__47471));
    InMux I__10997 (
            .O(N__47471),
            .I(N__47465));
    InMux I__10996 (
            .O(N__47470),
            .I(N__47465));
    LocalMux I__10995 (
            .O(N__47465),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__10994 (
            .O(N__47462),
            .I(N__47459));
    InMux I__10993 (
            .O(N__47459),
            .I(N__47456));
    LocalMux I__10992 (
            .O(N__47456),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt24 ));
    InMux I__10991 (
            .O(N__47453),
            .I(N__47449));
    InMux I__10990 (
            .O(N__47452),
            .I(N__47446));
    LocalMux I__10989 (
            .O(N__47449),
            .I(N__47440));
    LocalMux I__10988 (
            .O(N__47446),
            .I(N__47440));
    InMux I__10987 (
            .O(N__47445),
            .I(N__47437));
    Span4Mux_h I__10986 (
            .O(N__47440),
            .I(N__47434));
    LocalMux I__10985 (
            .O(N__47437),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__10984 (
            .O(N__47434),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    CascadeMux I__10983 (
            .O(N__47429),
            .I(N__47426));
    InMux I__10982 (
            .O(N__47426),
            .I(N__47422));
    InMux I__10981 (
            .O(N__47425),
            .I(N__47419));
    LocalMux I__10980 (
            .O(N__47422),
            .I(N__47413));
    LocalMux I__10979 (
            .O(N__47419),
            .I(N__47413));
    InMux I__10978 (
            .O(N__47418),
            .I(N__47410));
    Span4Mux_h I__10977 (
            .O(N__47413),
            .I(N__47407));
    LocalMux I__10976 (
            .O(N__47410),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__10975 (
            .O(N__47407),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__10974 (
            .O(N__47402),
            .I(N__47399));
    LocalMux I__10973 (
            .O(N__47399),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ));
    InMux I__10972 (
            .O(N__47396),
            .I(N__47393));
    LocalMux I__10971 (
            .O(N__47393),
            .I(N__47389));
    InMux I__10970 (
            .O(N__47392),
            .I(N__47386));
    Odrv12 I__10969 (
            .O(N__47389),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    LocalMux I__10968 (
            .O(N__47386),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    CascadeMux I__10967 (
            .O(N__47381),
            .I(elapsed_time_ns_1_RNI25DN9_0_24_cascade_));
    InMux I__10966 (
            .O(N__47378),
            .I(N__47373));
    InMux I__10965 (
            .O(N__47377),
            .I(N__47368));
    InMux I__10964 (
            .O(N__47376),
            .I(N__47368));
    LocalMux I__10963 (
            .O(N__47373),
            .I(N__47365));
    LocalMux I__10962 (
            .O(N__47368),
            .I(N__47362));
    Span4Mux_h I__10961 (
            .O(N__47365),
            .I(N__47357));
    Span4Mux_h I__10960 (
            .O(N__47362),
            .I(N__47357));
    Span4Mux_v I__10959 (
            .O(N__47357),
            .I(N__47353));
    InMux I__10958 (
            .O(N__47356),
            .I(N__47350));
    Odrv4 I__10957 (
            .O(N__47353),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__10956 (
            .O(N__47350),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__10955 (
            .O(N__47345),
            .I(N__47339));
    InMux I__10954 (
            .O(N__47344),
            .I(N__47339));
    LocalMux I__10953 (
            .O(N__47339),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    CascadeMux I__10952 (
            .O(N__47336),
            .I(N__47333));
    InMux I__10951 (
            .O(N__47333),
            .I(N__47330));
    LocalMux I__10950 (
            .O(N__47330),
            .I(N__47327));
    Span4Mux_h I__10949 (
            .O(N__47327),
            .I(N__47324));
    Span4Mux_h I__10948 (
            .O(N__47324),
            .I(N__47321));
    Odrv4 I__10947 (
            .O(N__47321),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__10946 (
            .O(N__47318),
            .I(N__47315));
    LocalMux I__10945 (
            .O(N__47315),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt20 ));
    InMux I__10944 (
            .O(N__47312),
            .I(N__47305));
    InMux I__10943 (
            .O(N__47311),
            .I(N__47305));
    InMux I__10942 (
            .O(N__47310),
            .I(N__47302));
    LocalMux I__10941 (
            .O(N__47305),
            .I(N__47299));
    LocalMux I__10940 (
            .O(N__47302),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__10939 (
            .O(N__47299),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    CascadeMux I__10938 (
            .O(N__47294),
            .I(N__47290));
    CascadeMux I__10937 (
            .O(N__47293),
            .I(N__47287));
    InMux I__10936 (
            .O(N__47290),
            .I(N__47281));
    InMux I__10935 (
            .O(N__47287),
            .I(N__47281));
    InMux I__10934 (
            .O(N__47286),
            .I(N__47278));
    LocalMux I__10933 (
            .O(N__47281),
            .I(N__47275));
    LocalMux I__10932 (
            .O(N__47278),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__10931 (
            .O(N__47275),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    CascadeMux I__10930 (
            .O(N__47270),
            .I(N__47267));
    InMux I__10929 (
            .O(N__47267),
            .I(N__47264));
    LocalMux I__10928 (
            .O(N__47264),
            .I(N__47261));
    Odrv4 I__10927 (
            .O(N__47261),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ));
    InMux I__10926 (
            .O(N__47258),
            .I(N__47255));
    LocalMux I__10925 (
            .O(N__47255),
            .I(N__47251));
    InMux I__10924 (
            .O(N__47254),
            .I(N__47247));
    Span4Mux_h I__10923 (
            .O(N__47251),
            .I(N__47244));
    InMux I__10922 (
            .O(N__47250),
            .I(N__47241));
    LocalMux I__10921 (
            .O(N__47247),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__10920 (
            .O(N__47244),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    LocalMux I__10919 (
            .O(N__47241),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__10918 (
            .O(N__47234),
            .I(N__47231));
    LocalMux I__10917 (
            .O(N__47231),
            .I(N__47228));
    Span4Mux_h I__10916 (
            .O(N__47228),
            .I(N__47222));
    InMux I__10915 (
            .O(N__47227),
            .I(N__47219));
    InMux I__10914 (
            .O(N__47226),
            .I(N__47214));
    InMux I__10913 (
            .O(N__47225),
            .I(N__47214));
    Odrv4 I__10912 (
            .O(N__47222),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__10911 (
            .O(N__47219),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__10910 (
            .O(N__47214),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    InMux I__10909 (
            .O(N__47207),
            .I(N__47204));
    LocalMux I__10908 (
            .O(N__47204),
            .I(N__47201));
    Span4Mux_h I__10907 (
            .O(N__47201),
            .I(N__47198));
    Odrv4 I__10906 (
            .O(N__47198),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__10905 (
            .O(N__47195),
            .I(N__47192));
    LocalMux I__10904 (
            .O(N__47192),
            .I(N__47187));
    InMux I__10903 (
            .O(N__47191),
            .I(N__47184));
    InMux I__10902 (
            .O(N__47190),
            .I(N__47181));
    Span4Mux_h I__10901 (
            .O(N__47187),
            .I(N__47178));
    LocalMux I__10900 (
            .O(N__47184),
            .I(N__47175));
    LocalMux I__10899 (
            .O(N__47181),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__10898 (
            .O(N__47178),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__10897 (
            .O(N__47175),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    CEMux I__10896 (
            .O(N__47168),
            .I(N__47144));
    CEMux I__10895 (
            .O(N__47167),
            .I(N__47144));
    CEMux I__10894 (
            .O(N__47166),
            .I(N__47144));
    CEMux I__10893 (
            .O(N__47165),
            .I(N__47144));
    CEMux I__10892 (
            .O(N__47164),
            .I(N__47144));
    CEMux I__10891 (
            .O(N__47163),
            .I(N__47144));
    CEMux I__10890 (
            .O(N__47162),
            .I(N__47144));
    CEMux I__10889 (
            .O(N__47161),
            .I(N__47144));
    GlobalMux I__10888 (
            .O(N__47144),
            .I(N__47141));
    gio2CtrlBuf I__10887 (
            .O(N__47141),
            .I(\current_shift_inst.timer_s1.N_167_i_g ));
    InMux I__10886 (
            .O(N__47138),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__10885 (
            .O(N__47135),
            .I(N__47131));
    InMux I__10884 (
            .O(N__47134),
            .I(N__47128));
    LocalMux I__10883 (
            .O(N__47131),
            .I(N__47125));
    LocalMux I__10882 (
            .O(N__47128),
            .I(N__47122));
    Span4Mux_v I__10881 (
            .O(N__47125),
            .I(N__47118));
    Span4Mux_h I__10880 (
            .O(N__47122),
            .I(N__47115));
    InMux I__10879 (
            .O(N__47121),
            .I(N__47112));
    Span4Mux_h I__10878 (
            .O(N__47118),
            .I(N__47109));
    Span4Mux_v I__10877 (
            .O(N__47115),
            .I(N__47106));
    LocalMux I__10876 (
            .O(N__47112),
            .I(N__47103));
    Odrv4 I__10875 (
            .O(N__47109),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__10874 (
            .O(N__47106),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__10873 (
            .O(N__47103),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__10872 (
            .O(N__47096),
            .I(N__47091));
    InMux I__10871 (
            .O(N__47095),
            .I(N__47087));
    InMux I__10870 (
            .O(N__47094),
            .I(N__47084));
    LocalMux I__10869 (
            .O(N__47091),
            .I(N__47081));
    InMux I__10868 (
            .O(N__47090),
            .I(N__47078));
    LocalMux I__10867 (
            .O(N__47087),
            .I(N__47075));
    LocalMux I__10866 (
            .O(N__47084),
            .I(N__47072));
    Span4Mux_h I__10865 (
            .O(N__47081),
            .I(N__47069));
    LocalMux I__10864 (
            .O(N__47078),
            .I(N__47066));
    Span4Mux_h I__10863 (
            .O(N__47075),
            .I(N__47063));
    Span4Mux_v I__10862 (
            .O(N__47072),
            .I(N__47060));
    Span4Mux_v I__10861 (
            .O(N__47069),
            .I(N__47053));
    Span4Mux_v I__10860 (
            .O(N__47066),
            .I(N__47053));
    Span4Mux_h I__10859 (
            .O(N__47063),
            .I(N__47053));
    Odrv4 I__10858 (
            .O(N__47060),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    Odrv4 I__10857 (
            .O(N__47053),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__10856 (
            .O(N__47048),
            .I(N__47045));
    LocalMux I__10855 (
            .O(N__47045),
            .I(N__47042));
    Span4Mux_v I__10854 (
            .O(N__47042),
            .I(N__47037));
    InMux I__10853 (
            .O(N__47041),
            .I(N__47034));
    InMux I__10852 (
            .O(N__47040),
            .I(N__47031));
    Span4Mux_v I__10851 (
            .O(N__47037),
            .I(N__47028));
    LocalMux I__10850 (
            .O(N__47034),
            .I(N__47025));
    LocalMux I__10849 (
            .O(N__47031),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    Odrv4 I__10848 (
            .O(N__47028),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    Odrv4 I__10847 (
            .O(N__47025),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    InMux I__10846 (
            .O(N__47018),
            .I(N__47015));
    LocalMux I__10845 (
            .O(N__47015),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    InMux I__10844 (
            .O(N__47012),
            .I(N__47009));
    LocalMux I__10843 (
            .O(N__47009),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    InMux I__10842 (
            .O(N__47006),
            .I(N__47003));
    LocalMux I__10841 (
            .O(N__47003),
            .I(N__47000));
    Span4Mux_v I__10840 (
            .O(N__47000),
            .I(N__46997));
    Span4Mux_h I__10839 (
            .O(N__46997),
            .I(N__46993));
    InMux I__10838 (
            .O(N__46996),
            .I(N__46990));
    Odrv4 I__10837 (
            .O(N__46993),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    LocalMux I__10836 (
            .O(N__46990),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    CascadeMux I__10835 (
            .O(N__46985),
            .I(elapsed_time_ns_1_RNI46CN9_0_17_cascade_));
    InMux I__10834 (
            .O(N__46982),
            .I(N__46976));
    InMux I__10833 (
            .O(N__46981),
            .I(N__46976));
    LocalMux I__10832 (
            .O(N__46976),
            .I(N__46972));
    InMux I__10831 (
            .O(N__46975),
            .I(N__46969));
    Span4Mux_h I__10830 (
            .O(N__46972),
            .I(N__46966));
    LocalMux I__10829 (
            .O(N__46969),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__10828 (
            .O(N__46966),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__10827 (
            .O(N__46961),
            .I(N__46957));
    CascadeMux I__10826 (
            .O(N__46960),
            .I(N__46954));
    InMux I__10825 (
            .O(N__46957),
            .I(N__46949));
    InMux I__10824 (
            .O(N__46954),
            .I(N__46949));
    LocalMux I__10823 (
            .O(N__46949),
            .I(N__46945));
    InMux I__10822 (
            .O(N__46948),
            .I(N__46942));
    Span4Mux_h I__10821 (
            .O(N__46945),
            .I(N__46939));
    LocalMux I__10820 (
            .O(N__46942),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__10819 (
            .O(N__46939),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__10818 (
            .O(N__46934),
            .I(N__46928));
    InMux I__10817 (
            .O(N__46933),
            .I(N__46928));
    LocalMux I__10816 (
            .O(N__46928),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__10815 (
            .O(N__46925),
            .I(N__46922));
    InMux I__10814 (
            .O(N__46922),
            .I(N__46919));
    LocalMux I__10813 (
            .O(N__46919),
            .I(N__46916));
    Odrv4 I__10812 (
            .O(N__46916),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    InMux I__10811 (
            .O(N__46913),
            .I(N__46910));
    LocalMux I__10810 (
            .O(N__46910),
            .I(N__46907));
    Span4Mux_v I__10809 (
            .O(N__46907),
            .I(N__46903));
    InMux I__10808 (
            .O(N__46906),
            .I(N__46900));
    Odrv4 I__10807 (
            .O(N__46903),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    LocalMux I__10806 (
            .O(N__46900),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    CascadeMux I__10805 (
            .O(N__46895),
            .I(elapsed_time_ns_1_RNI13CN9_0_14_cascade_));
    InMux I__10804 (
            .O(N__46892),
            .I(N__46889));
    LocalMux I__10803 (
            .O(N__46889),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__10802 (
            .O(N__46886),
            .I(N__46880));
    InMux I__10801 (
            .O(N__46885),
            .I(N__46880));
    LocalMux I__10800 (
            .O(N__46880),
            .I(N__46876));
    InMux I__10799 (
            .O(N__46879),
            .I(N__46873));
    Span4Mux_h I__10798 (
            .O(N__46876),
            .I(N__46870));
    LocalMux I__10797 (
            .O(N__46873),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__10796 (
            .O(N__46870),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    CascadeMux I__10795 (
            .O(N__46865),
            .I(N__46862));
    InMux I__10794 (
            .O(N__46862),
            .I(N__46858));
    InMux I__10793 (
            .O(N__46861),
            .I(N__46855));
    LocalMux I__10792 (
            .O(N__46858),
            .I(N__46851));
    LocalMux I__10791 (
            .O(N__46855),
            .I(N__46848));
    InMux I__10790 (
            .O(N__46854),
            .I(N__46845));
    Span4Mux_h I__10789 (
            .O(N__46851),
            .I(N__46840));
    Span4Mux_h I__10788 (
            .O(N__46848),
            .I(N__46840));
    LocalMux I__10787 (
            .O(N__46845),
            .I(N__46837));
    Span4Mux_v I__10786 (
            .O(N__46840),
            .I(N__46833));
    Span4Mux_h I__10785 (
            .O(N__46837),
            .I(N__46830));
    InMux I__10784 (
            .O(N__46836),
            .I(N__46827));
    Odrv4 I__10783 (
            .O(N__46833),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__10782 (
            .O(N__46830),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__10781 (
            .O(N__46827),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__10780 (
            .O(N__46820),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__10779 (
            .O(N__46817),
            .I(N__46811));
    InMux I__10778 (
            .O(N__46816),
            .I(N__46811));
    LocalMux I__10777 (
            .O(N__46811),
            .I(N__46807));
    InMux I__10776 (
            .O(N__46810),
            .I(N__46804));
    Span4Mux_h I__10775 (
            .O(N__46807),
            .I(N__46801));
    LocalMux I__10774 (
            .O(N__46804),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__10773 (
            .O(N__46801),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    CascadeMux I__10772 (
            .O(N__46796),
            .I(N__46792));
    InMux I__10771 (
            .O(N__46795),
            .I(N__46789));
    InMux I__10770 (
            .O(N__46792),
            .I(N__46786));
    LocalMux I__10769 (
            .O(N__46789),
            .I(N__46783));
    LocalMux I__10768 (
            .O(N__46786),
            .I(N__46779));
    Span4Mux_h I__10767 (
            .O(N__46783),
            .I(N__46776));
    InMux I__10766 (
            .O(N__46782),
            .I(N__46773));
    Span4Mux_h I__10765 (
            .O(N__46779),
            .I(N__46767));
    Span4Mux_v I__10764 (
            .O(N__46776),
            .I(N__46767));
    LocalMux I__10763 (
            .O(N__46773),
            .I(N__46764));
    InMux I__10762 (
            .O(N__46772),
            .I(N__46761));
    Odrv4 I__10761 (
            .O(N__46767),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__10760 (
            .O(N__46764),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__10759 (
            .O(N__46761),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__10758 (
            .O(N__46754),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__10757 (
            .O(N__46751),
            .I(N__46747));
    CascadeMux I__10756 (
            .O(N__46750),
            .I(N__46744));
    InMux I__10755 (
            .O(N__46747),
            .I(N__46739));
    InMux I__10754 (
            .O(N__46744),
            .I(N__46739));
    LocalMux I__10753 (
            .O(N__46739),
            .I(N__46735));
    InMux I__10752 (
            .O(N__46738),
            .I(N__46732));
    Span4Mux_h I__10751 (
            .O(N__46735),
            .I(N__46729));
    LocalMux I__10750 (
            .O(N__46732),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__10749 (
            .O(N__46729),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    CascadeMux I__10748 (
            .O(N__46724),
            .I(N__46721));
    InMux I__10747 (
            .O(N__46721),
            .I(N__46717));
    InMux I__10746 (
            .O(N__46720),
            .I(N__46713));
    LocalMux I__10745 (
            .O(N__46717),
            .I(N__46710));
    InMux I__10744 (
            .O(N__46716),
            .I(N__46707));
    LocalMux I__10743 (
            .O(N__46713),
            .I(N__46704));
    Span4Mux_v I__10742 (
            .O(N__46710),
            .I(N__46701));
    LocalMux I__10741 (
            .O(N__46707),
            .I(N__46698));
    Span4Mux_h I__10740 (
            .O(N__46704),
            .I(N__46694));
    Span4Mux_h I__10739 (
            .O(N__46701),
            .I(N__46691));
    Span12Mux_v I__10738 (
            .O(N__46698),
            .I(N__46688));
    InMux I__10737 (
            .O(N__46697),
            .I(N__46685));
    Odrv4 I__10736 (
            .O(N__46694),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__10735 (
            .O(N__46691),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv12 I__10734 (
            .O(N__46688),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__10733 (
            .O(N__46685),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__10732 (
            .O(N__46676),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__10731 (
            .O(N__46673),
            .I(N__46669));
    CascadeMux I__10730 (
            .O(N__46672),
            .I(N__46666));
    InMux I__10729 (
            .O(N__46669),
            .I(N__46661));
    InMux I__10728 (
            .O(N__46666),
            .I(N__46661));
    LocalMux I__10727 (
            .O(N__46661),
            .I(N__46657));
    InMux I__10726 (
            .O(N__46660),
            .I(N__46654));
    Span4Mux_h I__10725 (
            .O(N__46657),
            .I(N__46651));
    LocalMux I__10724 (
            .O(N__46654),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__10723 (
            .O(N__46651),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__10722 (
            .O(N__46646),
            .I(N__46642));
    InMux I__10721 (
            .O(N__46645),
            .I(N__46638));
    LocalMux I__10720 (
            .O(N__46642),
            .I(N__46635));
    InMux I__10719 (
            .O(N__46641),
            .I(N__46632));
    LocalMux I__10718 (
            .O(N__46638),
            .I(N__46629));
    Span4Mux_v I__10717 (
            .O(N__46635),
            .I(N__46624));
    LocalMux I__10716 (
            .O(N__46632),
            .I(N__46624));
    Span4Mux_h I__10715 (
            .O(N__46629),
            .I(N__46620));
    Span4Mux_h I__10714 (
            .O(N__46624),
            .I(N__46617));
    InMux I__10713 (
            .O(N__46623),
            .I(N__46614));
    Odrv4 I__10712 (
            .O(N__46620),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__10711 (
            .O(N__46617),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__10710 (
            .O(N__46614),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__10709 (
            .O(N__46607),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__10708 (
            .O(N__46604),
            .I(N__46601));
    InMux I__10707 (
            .O(N__46601),
            .I(N__46598));
    LocalMux I__10706 (
            .O(N__46598),
            .I(N__46594));
    InMux I__10705 (
            .O(N__46597),
            .I(N__46591));
    Span4Mux_v I__10704 (
            .O(N__46594),
            .I(N__46585));
    LocalMux I__10703 (
            .O(N__46591),
            .I(N__46585));
    InMux I__10702 (
            .O(N__46590),
            .I(N__46582));
    Span4Mux_h I__10701 (
            .O(N__46585),
            .I(N__46579));
    LocalMux I__10700 (
            .O(N__46582),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__10699 (
            .O(N__46579),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__10698 (
            .O(N__46574),
            .I(N__46571));
    LocalMux I__10697 (
            .O(N__46571),
            .I(N__46567));
    CascadeMux I__10696 (
            .O(N__46570),
            .I(N__46564));
    Span4Mux_h I__10695 (
            .O(N__46567),
            .I(N__46559));
    InMux I__10694 (
            .O(N__46564),
            .I(N__46554));
    InMux I__10693 (
            .O(N__46563),
            .I(N__46554));
    InMux I__10692 (
            .O(N__46562),
            .I(N__46551));
    Span4Mux_v I__10691 (
            .O(N__46559),
            .I(N__46544));
    LocalMux I__10690 (
            .O(N__46554),
            .I(N__46544));
    LocalMux I__10689 (
            .O(N__46551),
            .I(N__46544));
    Span4Mux_h I__10688 (
            .O(N__46544),
            .I(N__46541));
    Odrv4 I__10687 (
            .O(N__46541),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__10686 (
            .O(N__46538),
            .I(bfn_18_14_0_));
    CascadeMux I__10685 (
            .O(N__46535),
            .I(N__46532));
    InMux I__10684 (
            .O(N__46532),
            .I(N__46529));
    LocalMux I__10683 (
            .O(N__46529),
            .I(N__46525));
    InMux I__10682 (
            .O(N__46528),
            .I(N__46522));
    Span4Mux_v I__10681 (
            .O(N__46525),
            .I(N__46516));
    LocalMux I__10680 (
            .O(N__46522),
            .I(N__46516));
    InMux I__10679 (
            .O(N__46521),
            .I(N__46513));
    Span4Mux_h I__10678 (
            .O(N__46516),
            .I(N__46510));
    LocalMux I__10677 (
            .O(N__46513),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__10676 (
            .O(N__46510),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    CascadeMux I__10675 (
            .O(N__46505),
            .I(N__46502));
    InMux I__10674 (
            .O(N__46502),
            .I(N__46498));
    InMux I__10673 (
            .O(N__46501),
            .I(N__46494));
    LocalMux I__10672 (
            .O(N__46498),
            .I(N__46491));
    InMux I__10671 (
            .O(N__46497),
            .I(N__46488));
    LocalMux I__10670 (
            .O(N__46494),
            .I(N__46485));
    Span4Mux_h I__10669 (
            .O(N__46491),
            .I(N__46482));
    LocalMux I__10668 (
            .O(N__46488),
            .I(N__46479));
    Span4Mux_h I__10667 (
            .O(N__46485),
            .I(N__46475));
    Span4Mux_v I__10666 (
            .O(N__46482),
            .I(N__46472));
    Span4Mux_h I__10665 (
            .O(N__46479),
            .I(N__46469));
    InMux I__10664 (
            .O(N__46478),
            .I(N__46466));
    Odrv4 I__10663 (
            .O(N__46475),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__10662 (
            .O(N__46472),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__10661 (
            .O(N__46469),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__10660 (
            .O(N__46466),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__10659 (
            .O(N__46457),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__10658 (
            .O(N__46454),
            .I(N__46451));
    LocalMux I__10657 (
            .O(N__46451),
            .I(N__46447));
    InMux I__10656 (
            .O(N__46450),
            .I(N__46444));
    Span4Mux_h I__10655 (
            .O(N__46447),
            .I(N__46441));
    LocalMux I__10654 (
            .O(N__46444),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__10653 (
            .O(N__46441),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    CascadeMux I__10652 (
            .O(N__46436),
            .I(N__46433));
    InMux I__10651 (
            .O(N__46433),
            .I(N__46428));
    InMux I__10650 (
            .O(N__46432),
            .I(N__46425));
    InMux I__10649 (
            .O(N__46431),
            .I(N__46422));
    LocalMux I__10648 (
            .O(N__46428),
            .I(N__46417));
    LocalMux I__10647 (
            .O(N__46425),
            .I(N__46417));
    LocalMux I__10646 (
            .O(N__46422),
            .I(N__46412));
    Span4Mux_v I__10645 (
            .O(N__46417),
            .I(N__46412));
    Odrv4 I__10644 (
            .O(N__46412),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__10643 (
            .O(N__46409),
            .I(N__46403));
    InMux I__10642 (
            .O(N__46408),
            .I(N__46398));
    InMux I__10641 (
            .O(N__46407),
            .I(N__46398));
    InMux I__10640 (
            .O(N__46406),
            .I(N__46395));
    LocalMux I__10639 (
            .O(N__46403),
            .I(N__46392));
    LocalMux I__10638 (
            .O(N__46398),
            .I(N__46387));
    LocalMux I__10637 (
            .O(N__46395),
            .I(N__46387));
    Span4Mux_h I__10636 (
            .O(N__46392),
            .I(N__46384));
    Span4Mux_v I__10635 (
            .O(N__46387),
            .I(N__46381));
    Odrv4 I__10634 (
            .O(N__46384),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__10633 (
            .O(N__46381),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__10632 (
            .O(N__46376),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__10631 (
            .O(N__46373),
            .I(N__46370));
    LocalMux I__10630 (
            .O(N__46370),
            .I(N__46366));
    InMux I__10629 (
            .O(N__46369),
            .I(N__46363));
    Span4Mux_h I__10628 (
            .O(N__46366),
            .I(N__46360));
    LocalMux I__10627 (
            .O(N__46363),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__10626 (
            .O(N__46360),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CascadeMux I__10625 (
            .O(N__46355),
            .I(N__46352));
    InMux I__10624 (
            .O(N__46352),
            .I(N__46348));
    InMux I__10623 (
            .O(N__46351),
            .I(N__46345));
    LocalMux I__10622 (
            .O(N__46348),
            .I(N__46339));
    LocalMux I__10621 (
            .O(N__46345),
            .I(N__46339));
    InMux I__10620 (
            .O(N__46344),
            .I(N__46336));
    Span4Mux_v I__10619 (
            .O(N__46339),
            .I(N__46333));
    LocalMux I__10618 (
            .O(N__46336),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__10617 (
            .O(N__46333),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    CascadeMux I__10616 (
            .O(N__46328),
            .I(N__46325));
    InMux I__10615 (
            .O(N__46325),
            .I(N__46321));
    InMux I__10614 (
            .O(N__46324),
            .I(N__46317));
    LocalMux I__10613 (
            .O(N__46321),
            .I(N__46314));
    InMux I__10612 (
            .O(N__46320),
            .I(N__46311));
    LocalMux I__10611 (
            .O(N__46317),
            .I(N__46308));
    Span4Mux_v I__10610 (
            .O(N__46314),
            .I(N__46303));
    LocalMux I__10609 (
            .O(N__46311),
            .I(N__46303));
    Span4Mux_v I__10608 (
            .O(N__46308),
            .I(N__46299));
    Span4Mux_h I__10607 (
            .O(N__46303),
            .I(N__46296));
    InMux I__10606 (
            .O(N__46302),
            .I(N__46293));
    Odrv4 I__10605 (
            .O(N__46299),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__10604 (
            .O(N__46296),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__10603 (
            .O(N__46293),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__10602 (
            .O(N__46286),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    CascadeMux I__10601 (
            .O(N__46283),
            .I(N__46280));
    InMux I__10600 (
            .O(N__46280),
            .I(N__46276));
    InMux I__10599 (
            .O(N__46279),
            .I(N__46273));
    LocalMux I__10598 (
            .O(N__46276),
            .I(N__46267));
    LocalMux I__10597 (
            .O(N__46273),
            .I(N__46267));
    InMux I__10596 (
            .O(N__46272),
            .I(N__46264));
    Span4Mux_h I__10595 (
            .O(N__46267),
            .I(N__46261));
    LocalMux I__10594 (
            .O(N__46264),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__10593 (
            .O(N__46261),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    CascadeMux I__10592 (
            .O(N__46256),
            .I(N__46253));
    InMux I__10591 (
            .O(N__46253),
            .I(N__46249));
    InMux I__10590 (
            .O(N__46252),
            .I(N__46246));
    LocalMux I__10589 (
            .O(N__46249),
            .I(N__46242));
    LocalMux I__10588 (
            .O(N__46246),
            .I(N__46239));
    InMux I__10587 (
            .O(N__46245),
            .I(N__46236));
    Span4Mux_v I__10586 (
            .O(N__46242),
            .I(N__46229));
    Span4Mux_v I__10585 (
            .O(N__46239),
            .I(N__46229));
    LocalMux I__10584 (
            .O(N__46236),
            .I(N__46229));
    Span4Mux_h I__10583 (
            .O(N__46229),
            .I(N__46225));
    InMux I__10582 (
            .O(N__46228),
            .I(N__46222));
    Odrv4 I__10581 (
            .O(N__46225),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__10580 (
            .O(N__46222),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__10579 (
            .O(N__46217),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__10578 (
            .O(N__46214),
            .I(N__46208));
    InMux I__10577 (
            .O(N__46213),
            .I(N__46208));
    LocalMux I__10576 (
            .O(N__46208),
            .I(N__46204));
    InMux I__10575 (
            .O(N__46207),
            .I(N__46201));
    Span4Mux_h I__10574 (
            .O(N__46204),
            .I(N__46198));
    LocalMux I__10573 (
            .O(N__46201),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__10572 (
            .O(N__46198),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    CascadeMux I__10571 (
            .O(N__46193),
            .I(N__46190));
    InMux I__10570 (
            .O(N__46190),
            .I(N__46187));
    LocalMux I__10569 (
            .O(N__46187),
            .I(N__46184));
    Span4Mux_v I__10568 (
            .O(N__46184),
            .I(N__46180));
    InMux I__10567 (
            .O(N__46183),
            .I(N__46177));
    Span4Mux_h I__10566 (
            .O(N__46180),
            .I(N__46173));
    LocalMux I__10565 (
            .O(N__46177),
            .I(N__46170));
    InMux I__10564 (
            .O(N__46176),
            .I(N__46167));
    Span4Mux_h I__10563 (
            .O(N__46173),
            .I(N__46162));
    Span4Mux_h I__10562 (
            .O(N__46170),
            .I(N__46162));
    LocalMux I__10561 (
            .O(N__46167),
            .I(N__46159));
    Span4Mux_v I__10560 (
            .O(N__46162),
            .I(N__46155));
    Span4Mux_h I__10559 (
            .O(N__46159),
            .I(N__46152));
    InMux I__10558 (
            .O(N__46158),
            .I(N__46149));
    Odrv4 I__10557 (
            .O(N__46155),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__10556 (
            .O(N__46152),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__10555 (
            .O(N__46149),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__10554 (
            .O(N__46142),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__10553 (
            .O(N__46139),
            .I(N__46136));
    InMux I__10552 (
            .O(N__46136),
            .I(N__46132));
    InMux I__10551 (
            .O(N__46135),
            .I(N__46129));
    LocalMux I__10550 (
            .O(N__46132),
            .I(N__46123));
    LocalMux I__10549 (
            .O(N__46129),
            .I(N__46123));
    InMux I__10548 (
            .O(N__46128),
            .I(N__46120));
    Span4Mux_h I__10547 (
            .O(N__46123),
            .I(N__46117));
    LocalMux I__10546 (
            .O(N__46120),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__10545 (
            .O(N__46117),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    CascadeMux I__10544 (
            .O(N__46112),
            .I(N__46108));
    CascadeMux I__10543 (
            .O(N__46111),
            .I(N__46105));
    InMux I__10542 (
            .O(N__46108),
            .I(N__46102));
    InMux I__10541 (
            .O(N__46105),
            .I(N__46098));
    LocalMux I__10540 (
            .O(N__46102),
            .I(N__46095));
    InMux I__10539 (
            .O(N__46101),
            .I(N__46091));
    LocalMux I__10538 (
            .O(N__46098),
            .I(N__46088));
    Span4Mux_v I__10537 (
            .O(N__46095),
            .I(N__46085));
    InMux I__10536 (
            .O(N__46094),
            .I(N__46082));
    LocalMux I__10535 (
            .O(N__46091),
            .I(N__46079));
    Span4Mux_h I__10534 (
            .O(N__46088),
            .I(N__46072));
    Span4Mux_v I__10533 (
            .O(N__46085),
            .I(N__46072));
    LocalMux I__10532 (
            .O(N__46082),
            .I(N__46072));
    Odrv4 I__10531 (
            .O(N__46079),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__10530 (
            .O(N__46072),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__10529 (
            .O(N__46067),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__10528 (
            .O(N__46064),
            .I(N__46060));
    CascadeMux I__10527 (
            .O(N__46063),
            .I(N__46057));
    InMux I__10526 (
            .O(N__46060),
            .I(N__46052));
    InMux I__10525 (
            .O(N__46057),
            .I(N__46052));
    LocalMux I__10524 (
            .O(N__46052),
            .I(N__46048));
    InMux I__10523 (
            .O(N__46051),
            .I(N__46045));
    Span4Mux_h I__10522 (
            .O(N__46048),
            .I(N__46042));
    LocalMux I__10521 (
            .O(N__46045),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__10520 (
            .O(N__46042),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__10519 (
            .O(N__46037),
            .I(N__46032));
    InMux I__10518 (
            .O(N__46036),
            .I(N__46029));
    InMux I__10517 (
            .O(N__46035),
            .I(N__46025));
    LocalMux I__10516 (
            .O(N__46032),
            .I(N__46020));
    LocalMux I__10515 (
            .O(N__46029),
            .I(N__46020));
    InMux I__10514 (
            .O(N__46028),
            .I(N__46017));
    LocalMux I__10513 (
            .O(N__46025),
            .I(N__46014));
    Span4Mux_v I__10512 (
            .O(N__46020),
            .I(N__46009));
    LocalMux I__10511 (
            .O(N__46017),
            .I(N__46009));
    Odrv4 I__10510 (
            .O(N__46014),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__10509 (
            .O(N__46009),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__10508 (
            .O(N__46004),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__10507 (
            .O(N__46001),
            .I(N__45998));
    InMux I__10506 (
            .O(N__45998),
            .I(N__45995));
    LocalMux I__10505 (
            .O(N__45995),
            .I(N__45991));
    InMux I__10504 (
            .O(N__45994),
            .I(N__45988));
    Span4Mux_v I__10503 (
            .O(N__45991),
            .I(N__45982));
    LocalMux I__10502 (
            .O(N__45988),
            .I(N__45982));
    InMux I__10501 (
            .O(N__45987),
            .I(N__45979));
    Span4Mux_h I__10500 (
            .O(N__45982),
            .I(N__45976));
    LocalMux I__10499 (
            .O(N__45979),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__10498 (
            .O(N__45976),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    CascadeMux I__10497 (
            .O(N__45971),
            .I(N__45968));
    InMux I__10496 (
            .O(N__45968),
            .I(N__45964));
    InMux I__10495 (
            .O(N__45967),
            .I(N__45960));
    LocalMux I__10494 (
            .O(N__45964),
            .I(N__45957));
    InMux I__10493 (
            .O(N__45963),
            .I(N__45954));
    LocalMux I__10492 (
            .O(N__45960),
            .I(N__45951));
    Span4Mux_v I__10491 (
            .O(N__45957),
            .I(N__45946));
    LocalMux I__10490 (
            .O(N__45954),
            .I(N__45946));
    Span4Mux_v I__10489 (
            .O(N__45951),
            .I(N__45942));
    Span4Mux_v I__10488 (
            .O(N__45946),
            .I(N__45939));
    InMux I__10487 (
            .O(N__45945),
            .I(N__45936));
    Odrv4 I__10486 (
            .O(N__45942),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__10485 (
            .O(N__45939),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__10484 (
            .O(N__45936),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__10483 (
            .O(N__45929),
            .I(bfn_18_13_0_));
    CascadeMux I__10482 (
            .O(N__45926),
            .I(N__45923));
    InMux I__10481 (
            .O(N__45923),
            .I(N__45920));
    LocalMux I__10480 (
            .O(N__45920),
            .I(N__45916));
    InMux I__10479 (
            .O(N__45919),
            .I(N__45913));
    Span4Mux_v I__10478 (
            .O(N__45916),
            .I(N__45907));
    LocalMux I__10477 (
            .O(N__45913),
            .I(N__45907));
    InMux I__10476 (
            .O(N__45912),
            .I(N__45904));
    Span4Mux_h I__10475 (
            .O(N__45907),
            .I(N__45901));
    LocalMux I__10474 (
            .O(N__45904),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__10473 (
            .O(N__45901),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    CascadeMux I__10472 (
            .O(N__45896),
            .I(N__45892));
    InMux I__10471 (
            .O(N__45895),
            .I(N__45888));
    InMux I__10470 (
            .O(N__45892),
            .I(N__45885));
    CascadeMux I__10469 (
            .O(N__45891),
            .I(N__45882));
    LocalMux I__10468 (
            .O(N__45888),
            .I(N__45877));
    LocalMux I__10467 (
            .O(N__45885),
            .I(N__45877));
    InMux I__10466 (
            .O(N__45882),
            .I(N__45874));
    Span4Mux_h I__10465 (
            .O(N__45877),
            .I(N__45870));
    LocalMux I__10464 (
            .O(N__45874),
            .I(N__45867));
    InMux I__10463 (
            .O(N__45873),
            .I(N__45864));
    Odrv4 I__10462 (
            .O(N__45870),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__10461 (
            .O(N__45867),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__10460 (
            .O(N__45864),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__10459 (
            .O(N__45857),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__10458 (
            .O(N__45854),
            .I(N__45851));
    InMux I__10457 (
            .O(N__45851),
            .I(N__45847));
    InMux I__10456 (
            .O(N__45850),
            .I(N__45844));
    LocalMux I__10455 (
            .O(N__45847),
            .I(N__45838));
    LocalMux I__10454 (
            .O(N__45844),
            .I(N__45838));
    InMux I__10453 (
            .O(N__45843),
            .I(N__45835));
    Span4Mux_v I__10452 (
            .O(N__45838),
            .I(N__45832));
    LocalMux I__10451 (
            .O(N__45835),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__10450 (
            .O(N__45832),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    CascadeMux I__10449 (
            .O(N__45827),
            .I(N__45824));
    InMux I__10448 (
            .O(N__45824),
            .I(N__45820));
    InMux I__10447 (
            .O(N__45823),
            .I(N__45816));
    LocalMux I__10446 (
            .O(N__45820),
            .I(N__45813));
    InMux I__10445 (
            .O(N__45819),
            .I(N__45810));
    LocalMux I__10444 (
            .O(N__45816),
            .I(N__45807));
    Span4Mux_v I__10443 (
            .O(N__45813),
            .I(N__45804));
    LocalMux I__10442 (
            .O(N__45810),
            .I(N__45801));
    Span4Mux_v I__10441 (
            .O(N__45807),
            .I(N__45797));
    Span4Mux_v I__10440 (
            .O(N__45804),
            .I(N__45794));
    Span4Mux_h I__10439 (
            .O(N__45801),
            .I(N__45791));
    InMux I__10438 (
            .O(N__45800),
            .I(N__45788));
    Odrv4 I__10437 (
            .O(N__45797),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__10436 (
            .O(N__45794),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__10435 (
            .O(N__45791),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__10434 (
            .O(N__45788),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__10433 (
            .O(N__45779),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__10432 (
            .O(N__45776),
            .I(N__45773));
    InMux I__10431 (
            .O(N__45773),
            .I(N__45768));
    InMux I__10430 (
            .O(N__45772),
            .I(N__45765));
    InMux I__10429 (
            .O(N__45771),
            .I(N__45762));
    LocalMux I__10428 (
            .O(N__45768),
            .I(N__45757));
    LocalMux I__10427 (
            .O(N__45765),
            .I(N__45757));
    LocalMux I__10426 (
            .O(N__45762),
            .I(N__45752));
    Span4Mux_v I__10425 (
            .O(N__45757),
            .I(N__45752));
    Odrv4 I__10424 (
            .O(N__45752),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__10423 (
            .O(N__45749),
            .I(N__45740));
    InMux I__10422 (
            .O(N__45748),
            .I(N__45740));
    InMux I__10421 (
            .O(N__45747),
            .I(N__45740));
    LocalMux I__10420 (
            .O(N__45740),
            .I(N__45736));
    InMux I__10419 (
            .O(N__45739),
            .I(N__45733));
    Odrv4 I__10418 (
            .O(N__45736),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__10417 (
            .O(N__45733),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__10416 (
            .O(N__45728),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__10415 (
            .O(N__45725),
            .I(N__45722));
    InMux I__10414 (
            .O(N__45722),
            .I(N__45718));
    InMux I__10413 (
            .O(N__45721),
            .I(N__45715));
    LocalMux I__10412 (
            .O(N__45718),
            .I(N__45709));
    LocalMux I__10411 (
            .O(N__45715),
            .I(N__45709));
    InMux I__10410 (
            .O(N__45714),
            .I(N__45706));
    Span4Mux_h I__10409 (
            .O(N__45709),
            .I(N__45703));
    LocalMux I__10408 (
            .O(N__45706),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__10407 (
            .O(N__45703),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    CascadeMux I__10406 (
            .O(N__45698),
            .I(N__45695));
    InMux I__10405 (
            .O(N__45695),
            .I(N__45691));
    InMux I__10404 (
            .O(N__45694),
            .I(N__45688));
    LocalMux I__10403 (
            .O(N__45691),
            .I(N__45684));
    LocalMux I__10402 (
            .O(N__45688),
            .I(N__45681));
    InMux I__10401 (
            .O(N__45687),
            .I(N__45678));
    Span4Mux_h I__10400 (
            .O(N__45684),
            .I(N__45674));
    Span4Mux_v I__10399 (
            .O(N__45681),
            .I(N__45671));
    LocalMux I__10398 (
            .O(N__45678),
            .I(N__45668));
    InMux I__10397 (
            .O(N__45677),
            .I(N__45665));
    Span4Mux_v I__10396 (
            .O(N__45674),
            .I(N__45662));
    Span4Mux_h I__10395 (
            .O(N__45671),
            .I(N__45655));
    Span4Mux_v I__10394 (
            .O(N__45668),
            .I(N__45655));
    LocalMux I__10393 (
            .O(N__45665),
            .I(N__45655));
    Odrv4 I__10392 (
            .O(N__45662),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__10391 (
            .O(N__45655),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__10390 (
            .O(N__45650),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__10389 (
            .O(N__45647),
            .I(N__45641));
    InMux I__10388 (
            .O(N__45646),
            .I(N__45641));
    LocalMux I__10387 (
            .O(N__45641),
            .I(N__45637));
    InMux I__10386 (
            .O(N__45640),
            .I(N__45634));
    Span4Mux_h I__10385 (
            .O(N__45637),
            .I(N__45631));
    LocalMux I__10384 (
            .O(N__45634),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__10383 (
            .O(N__45631),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__10382 (
            .O(N__45626),
            .I(N__45623));
    LocalMux I__10381 (
            .O(N__45623),
            .I(N__45617));
    InMux I__10380 (
            .O(N__45622),
            .I(N__45612));
    InMux I__10379 (
            .O(N__45621),
            .I(N__45612));
    InMux I__10378 (
            .O(N__45620),
            .I(N__45609));
    Span4Mux_h I__10377 (
            .O(N__45617),
            .I(N__45606));
    LocalMux I__10376 (
            .O(N__45612),
            .I(N__45603));
    LocalMux I__10375 (
            .O(N__45609),
            .I(N__45600));
    Span4Mux_v I__10374 (
            .O(N__45606),
            .I(N__45597));
    Span4Mux_v I__10373 (
            .O(N__45603),
            .I(N__45592));
    Span4Mux_h I__10372 (
            .O(N__45600),
            .I(N__45592));
    Odrv4 I__10371 (
            .O(N__45597),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__10370 (
            .O(N__45592),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__10369 (
            .O(N__45587),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__10368 (
            .O(N__45584),
            .I(N__45578));
    InMux I__10367 (
            .O(N__45583),
            .I(N__45578));
    LocalMux I__10366 (
            .O(N__45578),
            .I(N__45574));
    InMux I__10365 (
            .O(N__45577),
            .I(N__45571));
    Span4Mux_h I__10364 (
            .O(N__45574),
            .I(N__45568));
    LocalMux I__10363 (
            .O(N__45571),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__10362 (
            .O(N__45568),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    CascadeMux I__10361 (
            .O(N__45563),
            .I(N__45559));
    CascadeMux I__10360 (
            .O(N__45562),
            .I(N__45556));
    InMux I__10359 (
            .O(N__45559),
            .I(N__45553));
    InMux I__10358 (
            .O(N__45556),
            .I(N__45550));
    LocalMux I__10357 (
            .O(N__45553),
            .I(N__45545));
    LocalMux I__10356 (
            .O(N__45550),
            .I(N__45542));
    InMux I__10355 (
            .O(N__45549),
            .I(N__45539));
    InMux I__10354 (
            .O(N__45548),
            .I(N__45536));
    Span4Mux_h I__10353 (
            .O(N__45545),
            .I(N__45531));
    Span4Mux_h I__10352 (
            .O(N__45542),
            .I(N__45531));
    LocalMux I__10351 (
            .O(N__45539),
            .I(N__45528));
    LocalMux I__10350 (
            .O(N__45536),
            .I(N__45525));
    Span4Mux_v I__10349 (
            .O(N__45531),
            .I(N__45522));
    Sp12to4 I__10348 (
            .O(N__45528),
            .I(N__45519));
    Span4Mux_h I__10347 (
            .O(N__45525),
            .I(N__45516));
    Odrv4 I__10346 (
            .O(N__45522),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv12 I__10345 (
            .O(N__45519),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__10344 (
            .O(N__45516),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__10343 (
            .O(N__45509),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__10342 (
            .O(N__45506),
            .I(N__45502));
    CascadeMux I__10341 (
            .O(N__45505),
            .I(N__45499));
    InMux I__10340 (
            .O(N__45502),
            .I(N__45494));
    InMux I__10339 (
            .O(N__45499),
            .I(N__45494));
    LocalMux I__10338 (
            .O(N__45494),
            .I(N__45490));
    InMux I__10337 (
            .O(N__45493),
            .I(N__45487));
    Span4Mux_h I__10336 (
            .O(N__45490),
            .I(N__45484));
    LocalMux I__10335 (
            .O(N__45487),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__10334 (
            .O(N__45484),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__10333 (
            .O(N__45479),
            .I(N__45471));
    InMux I__10332 (
            .O(N__45478),
            .I(N__45471));
    InMux I__10331 (
            .O(N__45477),
            .I(N__45468));
    InMux I__10330 (
            .O(N__45476),
            .I(N__45465));
    LocalMux I__10329 (
            .O(N__45471),
            .I(N__45462));
    LocalMux I__10328 (
            .O(N__45468),
            .I(N__45459));
    LocalMux I__10327 (
            .O(N__45465),
            .I(N__45454));
    Span4Mux_h I__10326 (
            .O(N__45462),
            .I(N__45454));
    Span12Mux_s10_v I__10325 (
            .O(N__45459),
            .I(N__45451));
    Span4Mux_h I__10324 (
            .O(N__45454),
            .I(N__45448));
    Odrv12 I__10323 (
            .O(N__45451),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv4 I__10322 (
            .O(N__45448),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__10321 (
            .O(N__45443),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__10320 (
            .O(N__45440),
            .I(N__45436));
    CascadeMux I__10319 (
            .O(N__45439),
            .I(N__45433));
    InMux I__10318 (
            .O(N__45436),
            .I(N__45430));
    InMux I__10317 (
            .O(N__45433),
            .I(N__45427));
    LocalMux I__10316 (
            .O(N__45430),
            .I(N__45423));
    LocalMux I__10315 (
            .O(N__45427),
            .I(N__45420));
    InMux I__10314 (
            .O(N__45426),
            .I(N__45417));
    Span4Mux_h I__10313 (
            .O(N__45423),
            .I(N__45414));
    Span4Mux_h I__10312 (
            .O(N__45420),
            .I(N__45411));
    LocalMux I__10311 (
            .O(N__45417),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__10310 (
            .O(N__45414),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__10309 (
            .O(N__45411),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    CascadeMux I__10308 (
            .O(N__45404),
            .I(N__45400));
    InMux I__10307 (
            .O(N__45403),
            .I(N__45397));
    InMux I__10306 (
            .O(N__45400),
            .I(N__45394));
    LocalMux I__10305 (
            .O(N__45397),
            .I(N__45390));
    LocalMux I__10304 (
            .O(N__45394),
            .I(N__45387));
    InMux I__10303 (
            .O(N__45393),
            .I(N__45384));
    Span4Mux_v I__10302 (
            .O(N__45390),
            .I(N__45379));
    Span4Mux_v I__10301 (
            .O(N__45387),
            .I(N__45379));
    LocalMux I__10300 (
            .O(N__45384),
            .I(N__45376));
    Span4Mux_h I__10299 (
            .O(N__45379),
            .I(N__45372));
    Span4Mux_h I__10298 (
            .O(N__45376),
            .I(N__45369));
    InMux I__10297 (
            .O(N__45375),
            .I(N__45366));
    Odrv4 I__10296 (
            .O(N__45372),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__10295 (
            .O(N__45369),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__10294 (
            .O(N__45366),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__10293 (
            .O(N__45359),
            .I(bfn_18_12_0_));
    CascadeMux I__10292 (
            .O(N__45356),
            .I(N__45353));
    InMux I__10291 (
            .O(N__45353),
            .I(N__45349));
    InMux I__10290 (
            .O(N__45352),
            .I(N__45346));
    LocalMux I__10289 (
            .O(N__45349),
            .I(N__45342));
    LocalMux I__10288 (
            .O(N__45346),
            .I(N__45339));
    InMux I__10287 (
            .O(N__45345),
            .I(N__45336));
    Span4Mux_h I__10286 (
            .O(N__45342),
            .I(N__45333));
    Span4Mux_h I__10285 (
            .O(N__45339),
            .I(N__45330));
    LocalMux I__10284 (
            .O(N__45336),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__10283 (
            .O(N__45333),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__10282 (
            .O(N__45330),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    CascadeMux I__10281 (
            .O(N__45323),
            .I(N__45319));
    InMux I__10280 (
            .O(N__45322),
            .I(N__45316));
    InMux I__10279 (
            .O(N__45319),
            .I(N__45313));
    LocalMux I__10278 (
            .O(N__45316),
            .I(N__45309));
    LocalMux I__10277 (
            .O(N__45313),
            .I(N__45306));
    InMux I__10276 (
            .O(N__45312),
            .I(N__45303));
    Span4Mux_h I__10275 (
            .O(N__45309),
            .I(N__45298));
    Span4Mux_h I__10274 (
            .O(N__45306),
            .I(N__45298));
    LocalMux I__10273 (
            .O(N__45303),
            .I(N__45295));
    Span4Mux_v I__10272 (
            .O(N__45298),
            .I(N__45291));
    Span4Mux_h I__10271 (
            .O(N__45295),
            .I(N__45288));
    InMux I__10270 (
            .O(N__45294),
            .I(N__45285));
    Odrv4 I__10269 (
            .O(N__45291),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__10268 (
            .O(N__45288),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__10267 (
            .O(N__45285),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__10266 (
            .O(N__45278),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__10265 (
            .O(N__45275),
            .I(N__45272));
    InMux I__10264 (
            .O(N__45272),
            .I(N__45268));
    InMux I__10263 (
            .O(N__45271),
            .I(N__45265));
    LocalMux I__10262 (
            .O(N__45268),
            .I(N__45259));
    LocalMux I__10261 (
            .O(N__45265),
            .I(N__45259));
    InMux I__10260 (
            .O(N__45264),
            .I(N__45256));
    Span4Mux_v I__10259 (
            .O(N__45259),
            .I(N__45253));
    LocalMux I__10258 (
            .O(N__45256),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__10257 (
            .O(N__45253),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    CascadeMux I__10256 (
            .O(N__45248),
            .I(N__45244));
    CascadeMux I__10255 (
            .O(N__45247),
            .I(N__45241));
    InMux I__10254 (
            .O(N__45244),
            .I(N__45238));
    InMux I__10253 (
            .O(N__45241),
            .I(N__45235));
    LocalMux I__10252 (
            .O(N__45238),
            .I(N__45232));
    LocalMux I__10251 (
            .O(N__45235),
            .I(N__45228));
    Span4Mux_v I__10250 (
            .O(N__45232),
            .I(N__45225));
    InMux I__10249 (
            .O(N__45231),
            .I(N__45222));
    Span4Mux_v I__10248 (
            .O(N__45228),
            .I(N__45218));
    Span4Mux_v I__10247 (
            .O(N__45225),
            .I(N__45215));
    LocalMux I__10246 (
            .O(N__45222),
            .I(N__45212));
    InMux I__10245 (
            .O(N__45221),
            .I(N__45209));
    Odrv4 I__10244 (
            .O(N__45218),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__10243 (
            .O(N__45215),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__10242 (
            .O(N__45212),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__10241 (
            .O(N__45209),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__10240 (
            .O(N__45200),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__10239 (
            .O(N__45197),
            .I(N__45194));
    InMux I__10238 (
            .O(N__45194),
            .I(N__45190));
    InMux I__10237 (
            .O(N__45193),
            .I(N__45187));
    LocalMux I__10236 (
            .O(N__45190),
            .I(N__45181));
    LocalMux I__10235 (
            .O(N__45187),
            .I(N__45181));
    InMux I__10234 (
            .O(N__45186),
            .I(N__45178));
    Span4Mux_v I__10233 (
            .O(N__45181),
            .I(N__45175));
    LocalMux I__10232 (
            .O(N__45178),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__10231 (
            .O(N__45175),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__10230 (
            .O(N__45170),
            .I(N__45166));
    CascadeMux I__10229 (
            .O(N__45169),
            .I(N__45163));
    LocalMux I__10228 (
            .O(N__45166),
            .I(N__45160));
    InMux I__10227 (
            .O(N__45163),
            .I(N__45157));
    Span4Mux_h I__10226 (
            .O(N__45160),
            .I(N__45152));
    LocalMux I__10225 (
            .O(N__45157),
            .I(N__45152));
    Span4Mux_v I__10224 (
            .O(N__45152),
            .I(N__45148));
    InMux I__10223 (
            .O(N__45151),
            .I(N__45145));
    Span4Mux_v I__10222 (
            .O(N__45148),
            .I(N__45141));
    LocalMux I__10221 (
            .O(N__45145),
            .I(N__45138));
    InMux I__10220 (
            .O(N__45144),
            .I(N__45135));
    Span4Mux_h I__10219 (
            .O(N__45141),
            .I(N__45132));
    Span4Mux_v I__10218 (
            .O(N__45138),
            .I(N__45127));
    LocalMux I__10217 (
            .O(N__45135),
            .I(N__45127));
    Odrv4 I__10216 (
            .O(N__45132),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__10215 (
            .O(N__45127),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__10214 (
            .O(N__45122),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__10213 (
            .O(N__45119),
            .I(N__45116));
    InMux I__10212 (
            .O(N__45116),
            .I(N__45113));
    LocalMux I__10211 (
            .O(N__45113),
            .I(N__45110));
    Odrv4 I__10210 (
            .O(N__45110),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__10209 (
            .O(N__45107),
            .I(N__45104));
    LocalMux I__10208 (
            .O(N__45104),
            .I(N__45101));
    Odrv4 I__10207 (
            .O(N__45101),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__10206 (
            .O(N__45098),
            .I(N__45084));
    CascadeMux I__10205 (
            .O(N__45097),
            .I(N__45080));
    CascadeMux I__10204 (
            .O(N__45096),
            .I(N__45076));
    CascadeMux I__10203 (
            .O(N__45095),
            .I(N__45072));
    CascadeMux I__10202 (
            .O(N__45094),
            .I(N__45068));
    CascadeMux I__10201 (
            .O(N__45093),
            .I(N__45064));
    CascadeMux I__10200 (
            .O(N__45092),
            .I(N__45060));
    CascadeMux I__10199 (
            .O(N__45091),
            .I(N__45055));
    CascadeMux I__10198 (
            .O(N__45090),
            .I(N__45051));
    CascadeMux I__10197 (
            .O(N__45089),
            .I(N__45047));
    InMux I__10196 (
            .O(N__45088),
            .I(N__45041));
    InMux I__10195 (
            .O(N__45087),
            .I(N__45021));
    InMux I__10194 (
            .O(N__45084),
            .I(N__45021));
    InMux I__10193 (
            .O(N__45083),
            .I(N__45021));
    InMux I__10192 (
            .O(N__45080),
            .I(N__45021));
    InMux I__10191 (
            .O(N__45079),
            .I(N__45021));
    InMux I__10190 (
            .O(N__45076),
            .I(N__45021));
    InMux I__10189 (
            .O(N__45075),
            .I(N__45021));
    InMux I__10188 (
            .O(N__45072),
            .I(N__45004));
    InMux I__10187 (
            .O(N__45071),
            .I(N__45004));
    InMux I__10186 (
            .O(N__45068),
            .I(N__45004));
    InMux I__10185 (
            .O(N__45067),
            .I(N__45004));
    InMux I__10184 (
            .O(N__45064),
            .I(N__45004));
    InMux I__10183 (
            .O(N__45063),
            .I(N__45004));
    InMux I__10182 (
            .O(N__45060),
            .I(N__45004));
    InMux I__10181 (
            .O(N__45059),
            .I(N__45004));
    InMux I__10180 (
            .O(N__45058),
            .I(N__44989));
    InMux I__10179 (
            .O(N__45055),
            .I(N__44989));
    InMux I__10178 (
            .O(N__45054),
            .I(N__44989));
    InMux I__10177 (
            .O(N__45051),
            .I(N__44989));
    InMux I__10176 (
            .O(N__45050),
            .I(N__44989));
    InMux I__10175 (
            .O(N__45047),
            .I(N__44989));
    InMux I__10174 (
            .O(N__45046),
            .I(N__44989));
    InMux I__10173 (
            .O(N__45045),
            .I(N__44978));
    InMux I__10172 (
            .O(N__45044),
            .I(N__44975));
    LocalMux I__10171 (
            .O(N__45041),
            .I(N__44972));
    InMux I__10170 (
            .O(N__45040),
            .I(N__44969));
    CascadeMux I__10169 (
            .O(N__45039),
            .I(N__44966));
    CascadeMux I__10168 (
            .O(N__45038),
            .I(N__44962));
    CascadeMux I__10167 (
            .O(N__45037),
            .I(N__44958));
    CascadeMux I__10166 (
            .O(N__45036),
            .I(N__44954));
    LocalMux I__10165 (
            .O(N__45021),
            .I(N__44950));
    LocalMux I__10164 (
            .O(N__45004),
            .I(N__44945));
    LocalMux I__10163 (
            .O(N__44989),
            .I(N__44945));
    InMux I__10162 (
            .O(N__44988),
            .I(N__44942));
    InMux I__10161 (
            .O(N__44987),
            .I(N__44935));
    InMux I__10160 (
            .O(N__44986),
            .I(N__44935));
    InMux I__10159 (
            .O(N__44985),
            .I(N__44935));
    InMux I__10158 (
            .O(N__44984),
            .I(N__44926));
    InMux I__10157 (
            .O(N__44983),
            .I(N__44926));
    InMux I__10156 (
            .O(N__44982),
            .I(N__44926));
    InMux I__10155 (
            .O(N__44981),
            .I(N__44926));
    LocalMux I__10154 (
            .O(N__44978),
            .I(N__44921));
    LocalMux I__10153 (
            .O(N__44975),
            .I(N__44914));
    Span4Mux_s1_v I__10152 (
            .O(N__44972),
            .I(N__44914));
    LocalMux I__10151 (
            .O(N__44969),
            .I(N__44914));
    InMux I__10150 (
            .O(N__44966),
            .I(N__44897));
    InMux I__10149 (
            .O(N__44965),
            .I(N__44897));
    InMux I__10148 (
            .O(N__44962),
            .I(N__44897));
    InMux I__10147 (
            .O(N__44961),
            .I(N__44897));
    InMux I__10146 (
            .O(N__44958),
            .I(N__44897));
    InMux I__10145 (
            .O(N__44957),
            .I(N__44897));
    InMux I__10144 (
            .O(N__44954),
            .I(N__44897));
    InMux I__10143 (
            .O(N__44953),
            .I(N__44897));
    Span4Mux_v I__10142 (
            .O(N__44950),
            .I(N__44892));
    Span4Mux_v I__10141 (
            .O(N__44945),
            .I(N__44892));
    LocalMux I__10140 (
            .O(N__44942),
            .I(N__44883));
    LocalMux I__10139 (
            .O(N__44935),
            .I(N__44883));
    LocalMux I__10138 (
            .O(N__44926),
            .I(N__44883));
    InMux I__10137 (
            .O(N__44925),
            .I(N__44880));
    CascadeMux I__10136 (
            .O(N__44924),
            .I(N__44869));
    Span12Mux_s5_v I__10135 (
            .O(N__44921),
            .I(N__44865));
    Span4Mux_h I__10134 (
            .O(N__44914),
            .I(N__44862));
    LocalMux I__10133 (
            .O(N__44897),
            .I(N__44859));
    Span4Mux_h I__10132 (
            .O(N__44892),
            .I(N__44856));
    InMux I__10131 (
            .O(N__44891),
            .I(N__44851));
    InMux I__10130 (
            .O(N__44890),
            .I(N__44851));
    Span4Mux_v I__10129 (
            .O(N__44883),
            .I(N__44848));
    LocalMux I__10128 (
            .O(N__44880),
            .I(N__44845));
    InMux I__10127 (
            .O(N__44879),
            .I(N__44838));
    InMux I__10126 (
            .O(N__44878),
            .I(N__44838));
    InMux I__10125 (
            .O(N__44877),
            .I(N__44838));
    InMux I__10124 (
            .O(N__44876),
            .I(N__44829));
    InMux I__10123 (
            .O(N__44875),
            .I(N__44829));
    InMux I__10122 (
            .O(N__44874),
            .I(N__44829));
    InMux I__10121 (
            .O(N__44873),
            .I(N__44829));
    InMux I__10120 (
            .O(N__44872),
            .I(N__44822));
    InMux I__10119 (
            .O(N__44869),
            .I(N__44822));
    InMux I__10118 (
            .O(N__44868),
            .I(N__44822));
    Span12Mux_v I__10117 (
            .O(N__44865),
            .I(N__44819));
    Sp12to4 I__10116 (
            .O(N__44862),
            .I(N__44816));
    Span12Mux_s9_h I__10115 (
            .O(N__44859),
            .I(N__44809));
    Sp12to4 I__10114 (
            .O(N__44856),
            .I(N__44809));
    LocalMux I__10113 (
            .O(N__44851),
            .I(N__44809));
    Span4Mux_v I__10112 (
            .O(N__44848),
            .I(N__44800));
    Span4Mux_v I__10111 (
            .O(N__44845),
            .I(N__44800));
    LocalMux I__10110 (
            .O(N__44838),
            .I(N__44800));
    LocalMux I__10109 (
            .O(N__44829),
            .I(N__44800));
    LocalMux I__10108 (
            .O(N__44822),
            .I(N__44797));
    Span12Mux_h I__10107 (
            .O(N__44819),
            .I(N__44794));
    Span12Mux_s10_v I__10106 (
            .O(N__44816),
            .I(N__44789));
    Span12Mux_h I__10105 (
            .O(N__44809),
            .I(N__44789));
    Span4Mux_h I__10104 (
            .O(N__44800),
            .I(N__44786));
    Span4Mux_v I__10103 (
            .O(N__44797),
            .I(N__44783));
    Odrv12 I__10102 (
            .O(N__44794),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__10101 (
            .O(N__44789),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__10100 (
            .O(N__44786),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__10099 (
            .O(N__44783),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__10098 (
            .O(N__44774),
            .I(N__44771));
    InMux I__10097 (
            .O(N__44771),
            .I(N__44768));
    LocalMux I__10096 (
            .O(N__44768),
            .I(N__44765));
    Span4Mux_v I__10095 (
            .O(N__44765),
            .I(N__44762));
    Odrv4 I__10094 (
            .O(N__44762),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__10093 (
            .O(N__44759),
            .I(N__44747));
    InMux I__10092 (
            .O(N__44758),
            .I(N__44747));
    InMux I__10091 (
            .O(N__44757),
            .I(N__44736));
    InMux I__10090 (
            .O(N__44756),
            .I(N__44736));
    InMux I__10089 (
            .O(N__44755),
            .I(N__44736));
    InMux I__10088 (
            .O(N__44754),
            .I(N__44736));
    InMux I__10087 (
            .O(N__44753),
            .I(N__44736));
    InMux I__10086 (
            .O(N__44752),
            .I(N__44701));
    LocalMux I__10085 (
            .O(N__44747),
            .I(N__44696));
    LocalMux I__10084 (
            .O(N__44736),
            .I(N__44696));
    InMux I__10083 (
            .O(N__44735),
            .I(N__44679));
    InMux I__10082 (
            .O(N__44734),
            .I(N__44679));
    InMux I__10081 (
            .O(N__44733),
            .I(N__44679));
    InMux I__10080 (
            .O(N__44732),
            .I(N__44679));
    InMux I__10079 (
            .O(N__44731),
            .I(N__44679));
    InMux I__10078 (
            .O(N__44730),
            .I(N__44679));
    InMux I__10077 (
            .O(N__44729),
            .I(N__44679));
    InMux I__10076 (
            .O(N__44728),
            .I(N__44679));
    InMux I__10075 (
            .O(N__44727),
            .I(N__44674));
    InMux I__10074 (
            .O(N__44726),
            .I(N__44669));
    InMux I__10073 (
            .O(N__44725),
            .I(N__44669));
    InMux I__10072 (
            .O(N__44724),
            .I(N__44642));
    InMux I__10071 (
            .O(N__44723),
            .I(N__44642));
    InMux I__10070 (
            .O(N__44722),
            .I(N__44642));
    InMux I__10069 (
            .O(N__44721),
            .I(N__44642));
    InMux I__10068 (
            .O(N__44720),
            .I(N__44642));
    InMux I__10067 (
            .O(N__44719),
            .I(N__44642));
    InMux I__10066 (
            .O(N__44718),
            .I(N__44642));
    InMux I__10065 (
            .O(N__44717),
            .I(N__44625));
    InMux I__10064 (
            .O(N__44716),
            .I(N__44625));
    InMux I__10063 (
            .O(N__44715),
            .I(N__44625));
    InMux I__10062 (
            .O(N__44714),
            .I(N__44625));
    InMux I__10061 (
            .O(N__44713),
            .I(N__44625));
    InMux I__10060 (
            .O(N__44712),
            .I(N__44625));
    InMux I__10059 (
            .O(N__44711),
            .I(N__44625));
    InMux I__10058 (
            .O(N__44710),
            .I(N__44625));
    InMux I__10057 (
            .O(N__44709),
            .I(N__44609));
    InMux I__10056 (
            .O(N__44708),
            .I(N__44609));
    InMux I__10055 (
            .O(N__44707),
            .I(N__44609));
    InMux I__10054 (
            .O(N__44706),
            .I(N__44609));
    InMux I__10053 (
            .O(N__44705),
            .I(N__44609));
    InMux I__10052 (
            .O(N__44704),
            .I(N__44606));
    LocalMux I__10051 (
            .O(N__44701),
            .I(N__44599));
    Span4Mux_h I__10050 (
            .O(N__44696),
            .I(N__44599));
    LocalMux I__10049 (
            .O(N__44679),
            .I(N__44599));
    InMux I__10048 (
            .O(N__44678),
            .I(N__44586));
    InMux I__10047 (
            .O(N__44677),
            .I(N__44586));
    LocalMux I__10046 (
            .O(N__44674),
            .I(N__44581));
    LocalMux I__10045 (
            .O(N__44669),
            .I(N__44581));
    InMux I__10044 (
            .O(N__44668),
            .I(N__44564));
    InMux I__10043 (
            .O(N__44667),
            .I(N__44564));
    InMux I__10042 (
            .O(N__44666),
            .I(N__44564));
    InMux I__10041 (
            .O(N__44665),
            .I(N__44564));
    InMux I__10040 (
            .O(N__44664),
            .I(N__44564));
    InMux I__10039 (
            .O(N__44663),
            .I(N__44564));
    InMux I__10038 (
            .O(N__44662),
            .I(N__44564));
    InMux I__10037 (
            .O(N__44661),
            .I(N__44564));
    InMux I__10036 (
            .O(N__44660),
            .I(N__44557));
    InMux I__10035 (
            .O(N__44659),
            .I(N__44557));
    InMux I__10034 (
            .O(N__44658),
            .I(N__44557));
    CascadeMux I__10033 (
            .O(N__44657),
            .I(N__44553));
    LocalMux I__10032 (
            .O(N__44642),
            .I(N__44545));
    LocalMux I__10031 (
            .O(N__44625),
            .I(N__44545));
    InMux I__10030 (
            .O(N__44624),
            .I(N__44534));
    InMux I__10029 (
            .O(N__44623),
            .I(N__44534));
    InMux I__10028 (
            .O(N__44622),
            .I(N__44534));
    InMux I__10027 (
            .O(N__44621),
            .I(N__44534));
    InMux I__10026 (
            .O(N__44620),
            .I(N__44534));
    LocalMux I__10025 (
            .O(N__44609),
            .I(N__44527));
    LocalMux I__10024 (
            .O(N__44606),
            .I(N__44527));
    Span4Mux_v I__10023 (
            .O(N__44599),
            .I(N__44527));
    InMux I__10022 (
            .O(N__44598),
            .I(N__44510));
    InMux I__10021 (
            .O(N__44597),
            .I(N__44510));
    InMux I__10020 (
            .O(N__44596),
            .I(N__44510));
    InMux I__10019 (
            .O(N__44595),
            .I(N__44510));
    InMux I__10018 (
            .O(N__44594),
            .I(N__44510));
    InMux I__10017 (
            .O(N__44593),
            .I(N__44510));
    InMux I__10016 (
            .O(N__44592),
            .I(N__44510));
    InMux I__10015 (
            .O(N__44591),
            .I(N__44510));
    LocalMux I__10014 (
            .O(N__44586),
            .I(N__44507));
    Span4Mux_h I__10013 (
            .O(N__44581),
            .I(N__44500));
    LocalMux I__10012 (
            .O(N__44564),
            .I(N__44500));
    LocalMux I__10011 (
            .O(N__44557),
            .I(N__44500));
    InMux I__10010 (
            .O(N__44556),
            .I(N__44489));
    InMux I__10009 (
            .O(N__44553),
            .I(N__44489));
    InMux I__10008 (
            .O(N__44552),
            .I(N__44489));
    InMux I__10007 (
            .O(N__44551),
            .I(N__44489));
    InMux I__10006 (
            .O(N__44550),
            .I(N__44489));
    Odrv12 I__10005 (
            .O(N__44545),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10004 (
            .O(N__44534),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10003 (
            .O(N__44527),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10002 (
            .O(N__44510),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10001 (
            .O(N__44507),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10000 (
            .O(N__44500),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__9999 (
            .O(N__44489),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__9998 (
            .O(N__44474),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__9997 (
            .O(N__44471),
            .I(N__44456));
    InMux I__9996 (
            .O(N__44470),
            .I(N__44456));
    InMux I__9995 (
            .O(N__44469),
            .I(N__44439));
    InMux I__9994 (
            .O(N__44468),
            .I(N__44439));
    InMux I__9993 (
            .O(N__44467),
            .I(N__44439));
    InMux I__9992 (
            .O(N__44466),
            .I(N__44439));
    InMux I__9991 (
            .O(N__44465),
            .I(N__44439));
    InMux I__9990 (
            .O(N__44464),
            .I(N__44439));
    InMux I__9989 (
            .O(N__44463),
            .I(N__44439));
    InMux I__9988 (
            .O(N__44462),
            .I(N__44439));
    InMux I__9987 (
            .O(N__44461),
            .I(N__44436));
    LocalMux I__9986 (
            .O(N__44456),
            .I(N__44433));
    LocalMux I__9985 (
            .O(N__44439),
            .I(N__44430));
    LocalMux I__9984 (
            .O(N__44436),
            .I(N__44421));
    Span4Mux_h I__9983 (
            .O(N__44433),
            .I(N__44421));
    Span4Mux_h I__9982 (
            .O(N__44430),
            .I(N__44418));
    InMux I__9981 (
            .O(N__44429),
            .I(N__44409));
    InMux I__9980 (
            .O(N__44428),
            .I(N__44409));
    InMux I__9979 (
            .O(N__44427),
            .I(N__44409));
    InMux I__9978 (
            .O(N__44426),
            .I(N__44409));
    Span4Mux_h I__9977 (
            .O(N__44421),
            .I(N__44406));
    Span4Mux_h I__9976 (
            .O(N__44418),
            .I(N__44403));
    LocalMux I__9975 (
            .O(N__44409),
            .I(N__44400));
    Odrv4 I__9974 (
            .O(N__44406),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__9973 (
            .O(N__44403),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv12 I__9972 (
            .O(N__44400),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__9971 (
            .O(N__44393),
            .I(N__44389));
    InMux I__9970 (
            .O(N__44392),
            .I(N__44386));
    LocalMux I__9969 (
            .O(N__44389),
            .I(N__44382));
    LocalMux I__9968 (
            .O(N__44386),
            .I(N__44379));
    InMux I__9967 (
            .O(N__44385),
            .I(N__44376));
    Span4Mux_v I__9966 (
            .O(N__44382),
            .I(N__44371));
    Span4Mux_h I__9965 (
            .O(N__44379),
            .I(N__44371));
    LocalMux I__9964 (
            .O(N__44376),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__9963 (
            .O(N__44371),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    CascadeMux I__9962 (
            .O(N__44366),
            .I(N__44363));
    InMux I__9961 (
            .O(N__44363),
            .I(N__44357));
    InMux I__9960 (
            .O(N__44362),
            .I(N__44357));
    LocalMux I__9959 (
            .O(N__44357),
            .I(N__44352));
    InMux I__9958 (
            .O(N__44356),
            .I(N__44349));
    InMux I__9957 (
            .O(N__44355),
            .I(N__44346));
    Span4Mux_h I__9956 (
            .O(N__44352),
            .I(N__44339));
    LocalMux I__9955 (
            .O(N__44349),
            .I(N__44339));
    LocalMux I__9954 (
            .O(N__44346),
            .I(N__44339));
    Odrv4 I__9953 (
            .O(N__44339),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__9952 (
            .O(N__44336),
            .I(N__44332));
    InMux I__9951 (
            .O(N__44335),
            .I(N__44329));
    LocalMux I__9950 (
            .O(N__44332),
            .I(N__44325));
    LocalMux I__9949 (
            .O(N__44329),
            .I(N__44322));
    InMux I__9948 (
            .O(N__44328),
            .I(N__44319));
    Span4Mux_h I__9947 (
            .O(N__44325),
            .I(N__44316));
    Odrv12 I__9946 (
            .O(N__44322),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__9945 (
            .O(N__44319),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__9944 (
            .O(N__44316),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    CascadeMux I__9943 (
            .O(N__44309),
            .I(N__44306));
    InMux I__9942 (
            .O(N__44306),
            .I(N__44302));
    InMux I__9941 (
            .O(N__44305),
            .I(N__44299));
    LocalMux I__9940 (
            .O(N__44302),
            .I(N__44295));
    LocalMux I__9939 (
            .O(N__44299),
            .I(N__44292));
    InMux I__9938 (
            .O(N__44298),
            .I(N__44289));
    Span4Mux_v I__9937 (
            .O(N__44295),
            .I(N__44285));
    Span4Mux_v I__9936 (
            .O(N__44292),
            .I(N__44280));
    LocalMux I__9935 (
            .O(N__44289),
            .I(N__44280));
    InMux I__9934 (
            .O(N__44288),
            .I(N__44277));
    Span4Mux_h I__9933 (
            .O(N__44285),
            .I(N__44274));
    Span4Mux_h I__9932 (
            .O(N__44280),
            .I(N__44269));
    LocalMux I__9931 (
            .O(N__44277),
            .I(N__44269));
    Odrv4 I__9930 (
            .O(N__44274),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__9929 (
            .O(N__44269),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__9928 (
            .O(N__44264),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__9927 (
            .O(N__44261),
            .I(N__44257));
    CascadeMux I__9926 (
            .O(N__44260),
            .I(N__44254));
    InMux I__9925 (
            .O(N__44257),
            .I(N__44249));
    InMux I__9924 (
            .O(N__44254),
            .I(N__44249));
    LocalMux I__9923 (
            .O(N__44249),
            .I(N__44245));
    InMux I__9922 (
            .O(N__44248),
            .I(N__44242));
    Span12Mux_s10_h I__9921 (
            .O(N__44245),
            .I(N__44239));
    LocalMux I__9920 (
            .O(N__44242),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__9919 (
            .O(N__44239),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    CascadeMux I__9918 (
            .O(N__44234),
            .I(N__44231));
    InMux I__9917 (
            .O(N__44231),
            .I(N__44227));
    InMux I__9916 (
            .O(N__44230),
            .I(N__44224));
    LocalMux I__9915 (
            .O(N__44227),
            .I(N__44219));
    LocalMux I__9914 (
            .O(N__44224),
            .I(N__44216));
    CascadeMux I__9913 (
            .O(N__44223),
            .I(N__44213));
    InMux I__9912 (
            .O(N__44222),
            .I(N__44210));
    Span4Mux_h I__9911 (
            .O(N__44219),
            .I(N__44205));
    Span4Mux_v I__9910 (
            .O(N__44216),
            .I(N__44205));
    InMux I__9909 (
            .O(N__44213),
            .I(N__44202));
    LocalMux I__9908 (
            .O(N__44210),
            .I(N__44199));
    Span4Mux_h I__9907 (
            .O(N__44205),
            .I(N__44196));
    LocalMux I__9906 (
            .O(N__44202),
            .I(N__44191));
    Span4Mux_h I__9905 (
            .O(N__44199),
            .I(N__44191));
    Odrv4 I__9904 (
            .O(N__44196),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__9903 (
            .O(N__44191),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__9902 (
            .O(N__44186),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__9901 (
            .O(N__44183),
            .I(N__44179));
    CascadeMux I__9900 (
            .O(N__44182),
            .I(N__44176));
    InMux I__9899 (
            .O(N__44179),
            .I(N__44171));
    InMux I__9898 (
            .O(N__44176),
            .I(N__44171));
    LocalMux I__9897 (
            .O(N__44171),
            .I(N__44167));
    InMux I__9896 (
            .O(N__44170),
            .I(N__44164));
    Span4Mux_v I__9895 (
            .O(N__44167),
            .I(N__44161));
    LocalMux I__9894 (
            .O(N__44164),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__9893 (
            .O(N__44161),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    CascadeMux I__9892 (
            .O(N__44156),
            .I(N__44152));
    CascadeMux I__9891 (
            .O(N__44155),
            .I(N__44149));
    InMux I__9890 (
            .O(N__44152),
            .I(N__44146));
    InMux I__9889 (
            .O(N__44149),
            .I(N__44143));
    LocalMux I__9888 (
            .O(N__44146),
            .I(N__44138));
    LocalMux I__9887 (
            .O(N__44143),
            .I(N__44138));
    Span4Mux_h I__9886 (
            .O(N__44138),
            .I(N__44133));
    InMux I__9885 (
            .O(N__44137),
            .I(N__44130));
    InMux I__9884 (
            .O(N__44136),
            .I(N__44127));
    Span4Mux_v I__9883 (
            .O(N__44133),
            .I(N__44124));
    LocalMux I__9882 (
            .O(N__44130),
            .I(N__44119));
    LocalMux I__9881 (
            .O(N__44127),
            .I(N__44119));
    Odrv4 I__9880 (
            .O(N__44124),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__9879 (
            .O(N__44119),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__9878 (
            .O(N__44114),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__9877 (
            .O(N__44111),
            .I(N__44108));
    InMux I__9876 (
            .O(N__44108),
            .I(N__44105));
    LocalMux I__9875 (
            .O(N__44105),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__9874 (
            .O(N__44102),
            .I(N__44099));
    LocalMux I__9873 (
            .O(N__44099),
            .I(N__44096));
    Odrv4 I__9872 (
            .O(N__44096),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__9871 (
            .O(N__44093),
            .I(N__44090));
    InMux I__9870 (
            .O(N__44090),
            .I(N__44087));
    LocalMux I__9869 (
            .O(N__44087),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__9868 (
            .O(N__44084),
            .I(N__44081));
    LocalMux I__9867 (
            .O(N__44081),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    CascadeMux I__9866 (
            .O(N__44078),
            .I(N__44075));
    InMux I__9865 (
            .O(N__44075),
            .I(N__44072));
    LocalMux I__9864 (
            .O(N__44072),
            .I(N__44069));
    Span12Mux_s9_h I__9863 (
            .O(N__44069),
            .I(N__44066));
    Odrv12 I__9862 (
            .O(N__44066),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__9861 (
            .O(N__44063),
            .I(N__44060));
    LocalMux I__9860 (
            .O(N__44060),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__9859 (
            .O(N__44057),
            .I(N__44054));
    InMux I__9858 (
            .O(N__44054),
            .I(N__44051));
    LocalMux I__9857 (
            .O(N__44051),
            .I(N__44048));
    Span4Mux_h I__9856 (
            .O(N__44048),
            .I(N__44045));
    Odrv4 I__9855 (
            .O(N__44045),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__9854 (
            .O(N__44042),
            .I(N__44039));
    LocalMux I__9853 (
            .O(N__44039),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    CascadeMux I__9852 (
            .O(N__44036),
            .I(N__44033));
    InMux I__9851 (
            .O(N__44033),
            .I(N__44030));
    LocalMux I__9850 (
            .O(N__44030),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__9849 (
            .O(N__44027),
            .I(N__44024));
    LocalMux I__9848 (
            .O(N__44024),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__9847 (
            .O(N__44021),
            .I(N__44018));
    InMux I__9846 (
            .O(N__44018),
            .I(N__44015));
    LocalMux I__9845 (
            .O(N__44015),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__9844 (
            .O(N__44012),
            .I(N__44009));
    LocalMux I__9843 (
            .O(N__44009),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__9842 (
            .O(N__44006),
            .I(N__44003));
    InMux I__9841 (
            .O(N__44003),
            .I(N__44000));
    LocalMux I__9840 (
            .O(N__44000),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    InMux I__9839 (
            .O(N__43997),
            .I(N__43994));
    LocalMux I__9838 (
            .O(N__43994),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__9837 (
            .O(N__43991),
            .I(N__43988));
    InMux I__9836 (
            .O(N__43988),
            .I(N__43985));
    LocalMux I__9835 (
            .O(N__43985),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__9834 (
            .O(N__43982),
            .I(N__43979));
    LocalMux I__9833 (
            .O(N__43979),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    CascadeMux I__9832 (
            .O(N__43976),
            .I(N__43973));
    InMux I__9831 (
            .O(N__43973),
            .I(N__43970));
    LocalMux I__9830 (
            .O(N__43970),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__9829 (
            .O(N__43967),
            .I(N__43964));
    LocalMux I__9828 (
            .O(N__43964),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__9827 (
            .O(N__43961),
            .I(N__43958));
    InMux I__9826 (
            .O(N__43958),
            .I(N__43955));
    LocalMux I__9825 (
            .O(N__43955),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__9824 (
            .O(N__43952),
            .I(N__43949));
    LocalMux I__9823 (
            .O(N__43949),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__9822 (
            .O(N__43946),
            .I(N__43943));
    InMux I__9821 (
            .O(N__43943),
            .I(N__43940));
    LocalMux I__9820 (
            .O(N__43940),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__9819 (
            .O(N__43937),
            .I(N__43934));
    InMux I__9818 (
            .O(N__43934),
            .I(N__43931));
    LocalMux I__9817 (
            .O(N__43931),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__9816 (
            .O(N__43928),
            .I(N__43925));
    LocalMux I__9815 (
            .O(N__43925),
            .I(N__43922));
    Span4Mux_h I__9814 (
            .O(N__43922),
            .I(N__43919));
    Span4Mux_h I__9813 (
            .O(N__43919),
            .I(N__43916));
    Odrv4 I__9812 (
            .O(N__43916),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__9811 (
            .O(N__43913),
            .I(N__43910));
    InMux I__9810 (
            .O(N__43910),
            .I(N__43907));
    LocalMux I__9809 (
            .O(N__43907),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__9808 (
            .O(N__43904),
            .I(N__43901));
    LocalMux I__9807 (
            .O(N__43901),
            .I(N__43898));
    Odrv12 I__9806 (
            .O(N__43898),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__9805 (
            .O(N__43895),
            .I(N__43889));
    InMux I__9804 (
            .O(N__43894),
            .I(N__43884));
    InMux I__9803 (
            .O(N__43893),
            .I(N__43884));
    InMux I__9802 (
            .O(N__43892),
            .I(N__43881));
    LocalMux I__9801 (
            .O(N__43889),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__9800 (
            .O(N__43884),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__9799 (
            .O(N__43881),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__9798 (
            .O(N__43874),
            .I(N__43870));
    InMux I__9797 (
            .O(N__43873),
            .I(N__43867));
    LocalMux I__9796 (
            .O(N__43870),
            .I(N__43863));
    LocalMux I__9795 (
            .O(N__43867),
            .I(N__43859));
    InMux I__9794 (
            .O(N__43866),
            .I(N__43856));
    Span4Mux_h I__9793 (
            .O(N__43863),
            .I(N__43853));
    InMux I__9792 (
            .O(N__43862),
            .I(N__43850));
    Odrv12 I__9791 (
            .O(N__43859),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    LocalMux I__9790 (
            .O(N__43856),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__9789 (
            .O(N__43853),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    LocalMux I__9788 (
            .O(N__43850),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__9787 (
            .O(N__43841),
            .I(N__43837));
    InMux I__9786 (
            .O(N__43840),
            .I(N__43833));
    LocalMux I__9785 (
            .O(N__43837),
            .I(N__43830));
    InMux I__9784 (
            .O(N__43836),
            .I(N__43827));
    LocalMux I__9783 (
            .O(N__43833),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    Odrv12 I__9782 (
            .O(N__43830),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__9781 (
            .O(N__43827),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    InMux I__9780 (
            .O(N__43820),
            .I(N__43817));
    LocalMux I__9779 (
            .O(N__43817),
            .I(N__43814));
    Span12Mux_v I__9778 (
            .O(N__43814),
            .I(N__43811));
    Odrv12 I__9777 (
            .O(N__43811),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__9776 (
            .O(N__43808),
            .I(N__43804));
    InMux I__9775 (
            .O(N__43807),
            .I(N__43801));
    LocalMux I__9774 (
            .O(N__43804),
            .I(N__43795));
    LocalMux I__9773 (
            .O(N__43801),
            .I(N__43792));
    InMux I__9772 (
            .O(N__43800),
            .I(N__43789));
    InMux I__9771 (
            .O(N__43799),
            .I(N__43784));
    InMux I__9770 (
            .O(N__43798),
            .I(N__43784));
    Span4Mux_h I__9769 (
            .O(N__43795),
            .I(N__43781));
    Odrv12 I__9768 (
            .O(N__43792),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__9767 (
            .O(N__43789),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__9766 (
            .O(N__43784),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__9765 (
            .O(N__43781),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__9764 (
            .O(N__43772),
            .I(N__43769));
    InMux I__9763 (
            .O(N__43769),
            .I(N__43766));
    LocalMux I__9762 (
            .O(N__43766),
            .I(N__43762));
    InMux I__9761 (
            .O(N__43765),
            .I(N__43759));
    Span4Mux_h I__9760 (
            .O(N__43762),
            .I(N__43756));
    LocalMux I__9759 (
            .O(N__43759),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv4 I__9758 (
            .O(N__43756),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    CascadeMux I__9757 (
            .O(N__43751),
            .I(N__43748));
    InMux I__9756 (
            .O(N__43748),
            .I(N__43745));
    LocalMux I__9755 (
            .O(N__43745),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__9754 (
            .O(N__43742),
            .I(N__43739));
    LocalMux I__9753 (
            .O(N__43739),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__9752 (
            .O(N__43736),
            .I(N__43731));
    CascadeMux I__9751 (
            .O(N__43735),
            .I(N__43728));
    InMux I__9750 (
            .O(N__43734),
            .I(N__43720));
    InMux I__9749 (
            .O(N__43731),
            .I(N__43720));
    InMux I__9748 (
            .O(N__43728),
            .I(N__43720));
    InMux I__9747 (
            .O(N__43727),
            .I(N__43717));
    LocalMux I__9746 (
            .O(N__43720),
            .I(N__43714));
    LocalMux I__9745 (
            .O(N__43717),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__9744 (
            .O(N__43714),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__9743 (
            .O(N__43709),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__9742 (
            .O(N__43706),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    CascadeMux I__9741 (
            .O(N__43703),
            .I(N__43700));
    InMux I__9740 (
            .O(N__43700),
            .I(N__43691));
    InMux I__9739 (
            .O(N__43699),
            .I(N__43691));
    InMux I__9738 (
            .O(N__43698),
            .I(N__43691));
    LocalMux I__9737 (
            .O(N__43691),
            .I(N__43687));
    InMux I__9736 (
            .O(N__43690),
            .I(N__43684));
    Span4Mux_h I__9735 (
            .O(N__43687),
            .I(N__43681));
    LocalMux I__9734 (
            .O(N__43684),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__9733 (
            .O(N__43681),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__9732 (
            .O(N__43676),
            .I(N__43673));
    InMux I__9731 (
            .O(N__43673),
            .I(N__43670));
    LocalMux I__9730 (
            .O(N__43670),
            .I(N__43667));
    Span4Mux_v I__9729 (
            .O(N__43667),
            .I(N__43664));
    Odrv4 I__9728 (
            .O(N__43664),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt28 ));
    InMux I__9727 (
            .O(N__43661),
            .I(N__43656));
    InMux I__9726 (
            .O(N__43660),
            .I(N__43651));
    InMux I__9725 (
            .O(N__43659),
            .I(N__43651));
    LocalMux I__9724 (
            .O(N__43656),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__9723 (
            .O(N__43651),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    CascadeMux I__9722 (
            .O(N__43646),
            .I(N__43643));
    InMux I__9721 (
            .O(N__43643),
            .I(N__43636));
    InMux I__9720 (
            .O(N__43642),
            .I(N__43636));
    InMux I__9719 (
            .O(N__43641),
            .I(N__43633));
    LocalMux I__9718 (
            .O(N__43636),
            .I(N__43630));
    LocalMux I__9717 (
            .O(N__43633),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__9716 (
            .O(N__43630),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__9715 (
            .O(N__43625),
            .I(N__43622));
    LocalMux I__9714 (
            .O(N__43622),
            .I(N__43619));
    Odrv12 I__9713 (
            .O(N__43619),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ));
    InMux I__9712 (
            .O(N__43616),
            .I(N__43613));
    LocalMux I__9711 (
            .O(N__43613),
            .I(N__43609));
    InMux I__9710 (
            .O(N__43612),
            .I(N__43606));
    Odrv4 I__9709 (
            .O(N__43609),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    LocalMux I__9708 (
            .O(N__43606),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    CascadeMux I__9707 (
            .O(N__43601),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_));
    CascadeMux I__9706 (
            .O(N__43598),
            .I(N__43595));
    InMux I__9705 (
            .O(N__43595),
            .I(N__43589));
    InMux I__9704 (
            .O(N__43594),
            .I(N__43589));
    LocalMux I__9703 (
            .O(N__43589),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    InMux I__9702 (
            .O(N__43586),
            .I(N__43580));
    InMux I__9701 (
            .O(N__43585),
            .I(N__43577));
    InMux I__9700 (
            .O(N__43584),
            .I(N__43574));
    InMux I__9699 (
            .O(N__43583),
            .I(N__43571));
    LocalMux I__9698 (
            .O(N__43580),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    LocalMux I__9697 (
            .O(N__43577),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    LocalMux I__9696 (
            .O(N__43574),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    LocalMux I__9695 (
            .O(N__43571),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__9694 (
            .O(N__43562),
            .I(N__43559));
    LocalMux I__9693 (
            .O(N__43559),
            .I(N__43555));
    InMux I__9692 (
            .O(N__43558),
            .I(N__43551));
    Span4Mux_h I__9691 (
            .O(N__43555),
            .I(N__43548));
    InMux I__9690 (
            .O(N__43554),
            .I(N__43545));
    LocalMux I__9689 (
            .O(N__43551),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    Odrv4 I__9688 (
            .O(N__43548),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    LocalMux I__9687 (
            .O(N__43545),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    InMux I__9686 (
            .O(N__43538),
            .I(N__43532));
    InMux I__9685 (
            .O(N__43537),
            .I(N__43532));
    LocalMux I__9684 (
            .O(N__43532),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    InMux I__9683 (
            .O(N__43529),
            .I(N__43526));
    LocalMux I__9682 (
            .O(N__43526),
            .I(N__43521));
    InMux I__9681 (
            .O(N__43525),
            .I(N__43516));
    InMux I__9680 (
            .O(N__43524),
            .I(N__43516));
    Span4Mux_h I__9679 (
            .O(N__43521),
            .I(N__43512));
    LocalMux I__9678 (
            .O(N__43516),
            .I(N__43509));
    InMux I__9677 (
            .O(N__43515),
            .I(N__43506));
    Odrv4 I__9676 (
            .O(N__43512),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv12 I__9675 (
            .O(N__43509),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__9674 (
            .O(N__43506),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__9673 (
            .O(N__43499),
            .I(N__43494));
    InMux I__9672 (
            .O(N__43498),
            .I(N__43489));
    InMux I__9671 (
            .O(N__43497),
            .I(N__43489));
    LocalMux I__9670 (
            .O(N__43494),
            .I(N__43486));
    LocalMux I__9669 (
            .O(N__43489),
            .I(N__43483));
    Span4Mux_v I__9668 (
            .O(N__43486),
            .I(N__43479));
    Span4Mux_v I__9667 (
            .O(N__43483),
            .I(N__43476));
    InMux I__9666 (
            .O(N__43482),
            .I(N__43473));
    Odrv4 I__9665 (
            .O(N__43479),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    Odrv4 I__9664 (
            .O(N__43476),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__9663 (
            .O(N__43473),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__9662 (
            .O(N__43466),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__9661 (
            .O(N__43463),
            .I(N__43458));
    InMux I__9660 (
            .O(N__43462),
            .I(N__43455));
    InMux I__9659 (
            .O(N__43461),
            .I(N__43450));
    InMux I__9658 (
            .O(N__43458),
            .I(N__43450));
    LocalMux I__9657 (
            .O(N__43455),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    LocalMux I__9656 (
            .O(N__43450),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__9655 (
            .O(N__43445),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    CascadeMux I__9654 (
            .O(N__43442),
            .I(N__43437));
    InMux I__9653 (
            .O(N__43441),
            .I(N__43434));
    InMux I__9652 (
            .O(N__43440),
            .I(N__43429));
    InMux I__9651 (
            .O(N__43437),
            .I(N__43429));
    LocalMux I__9650 (
            .O(N__43434),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    LocalMux I__9649 (
            .O(N__43429),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__9648 (
            .O(N__43424),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__9647 (
            .O(N__43421),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__9646 (
            .O(N__43418),
            .I(bfn_17_21_0_));
    InMux I__9645 (
            .O(N__43415),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__9644 (
            .O(N__43412),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__9643 (
            .O(N__43409),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__9642 (
            .O(N__43406),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__9641 (
            .O(N__43403),
            .I(N__43399));
    InMux I__9640 (
            .O(N__43402),
            .I(N__43396));
    LocalMux I__9639 (
            .O(N__43399),
            .I(N__43393));
    LocalMux I__9638 (
            .O(N__43396),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__9637 (
            .O(N__43393),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__9636 (
            .O(N__43388),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__9635 (
            .O(N__43385),
            .I(N__43381));
    InMux I__9634 (
            .O(N__43384),
            .I(N__43378));
    LocalMux I__9633 (
            .O(N__43381),
            .I(N__43375));
    LocalMux I__9632 (
            .O(N__43378),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__9631 (
            .O(N__43375),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__9630 (
            .O(N__43370),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__9629 (
            .O(N__43367),
            .I(N__43363));
    InMux I__9628 (
            .O(N__43366),
            .I(N__43360));
    LocalMux I__9627 (
            .O(N__43363),
            .I(N__43357));
    LocalMux I__9626 (
            .O(N__43360),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__9625 (
            .O(N__43357),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__9624 (
            .O(N__43352),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__9623 (
            .O(N__43349),
            .I(N__43346));
    LocalMux I__9622 (
            .O(N__43346),
            .I(N__43342));
    InMux I__9621 (
            .O(N__43345),
            .I(N__43339));
    Span4Mux_v I__9620 (
            .O(N__43342),
            .I(N__43336));
    LocalMux I__9619 (
            .O(N__43339),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__9618 (
            .O(N__43336),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__9617 (
            .O(N__43331),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__9616 (
            .O(N__43328),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__9615 (
            .O(N__43325),
            .I(bfn_17_20_0_));
    InMux I__9614 (
            .O(N__43322),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__9613 (
            .O(N__43319),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__9612 (
            .O(N__43316),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__9611 (
            .O(N__43313),
            .I(N__43309));
    InMux I__9610 (
            .O(N__43312),
            .I(N__43306));
    LocalMux I__9609 (
            .O(N__43309),
            .I(N__43303));
    LocalMux I__9608 (
            .O(N__43306),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__9607 (
            .O(N__43303),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__9606 (
            .O(N__43298),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__9605 (
            .O(N__43295),
            .I(N__43291));
    InMux I__9604 (
            .O(N__43294),
            .I(N__43288));
    LocalMux I__9603 (
            .O(N__43291),
            .I(N__43285));
    LocalMux I__9602 (
            .O(N__43288),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__9601 (
            .O(N__43285),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__9600 (
            .O(N__43280),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__9599 (
            .O(N__43277),
            .I(N__43273));
    InMux I__9598 (
            .O(N__43276),
            .I(N__43270));
    LocalMux I__9597 (
            .O(N__43273),
            .I(N__43267));
    LocalMux I__9596 (
            .O(N__43270),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__9595 (
            .O(N__43267),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__9594 (
            .O(N__43262),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__9593 (
            .O(N__43259),
            .I(N__43255));
    InMux I__9592 (
            .O(N__43258),
            .I(N__43252));
    LocalMux I__9591 (
            .O(N__43255),
            .I(N__43249));
    LocalMux I__9590 (
            .O(N__43252),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv12 I__9589 (
            .O(N__43249),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__9588 (
            .O(N__43244),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__9587 (
            .O(N__43241),
            .I(N__43237));
    InMux I__9586 (
            .O(N__43240),
            .I(N__43234));
    LocalMux I__9585 (
            .O(N__43237),
            .I(N__43231));
    LocalMux I__9584 (
            .O(N__43234),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv12 I__9583 (
            .O(N__43231),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__9582 (
            .O(N__43226),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__9581 (
            .O(N__43223),
            .I(N__43219));
    InMux I__9580 (
            .O(N__43222),
            .I(N__43216));
    LocalMux I__9579 (
            .O(N__43219),
            .I(N__43213));
    LocalMux I__9578 (
            .O(N__43216),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__9577 (
            .O(N__43213),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__9576 (
            .O(N__43208),
            .I(bfn_17_19_0_));
    InMux I__9575 (
            .O(N__43205),
            .I(N__43202));
    LocalMux I__9574 (
            .O(N__43202),
            .I(N__43198));
    InMux I__9573 (
            .O(N__43201),
            .I(N__43195));
    Span4Mux_h I__9572 (
            .O(N__43198),
            .I(N__43192));
    LocalMux I__9571 (
            .O(N__43195),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__9570 (
            .O(N__43192),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__9569 (
            .O(N__43187),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__9568 (
            .O(N__43184),
            .I(N__43180));
    InMux I__9567 (
            .O(N__43183),
            .I(N__43177));
    LocalMux I__9566 (
            .O(N__43180),
            .I(N__43174));
    LocalMux I__9565 (
            .O(N__43177),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__9564 (
            .O(N__43174),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__9563 (
            .O(N__43169),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__9562 (
            .O(N__43166),
            .I(N__43163));
    LocalMux I__9561 (
            .O(N__43163),
            .I(N__43160));
    Span4Mux_h I__9560 (
            .O(N__43160),
            .I(N__43157));
    Odrv4 I__9559 (
            .O(N__43157),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ));
    CascadeMux I__9558 (
            .O(N__43154),
            .I(N__43151));
    InMux I__9557 (
            .O(N__43151),
            .I(N__43148));
    LocalMux I__9556 (
            .O(N__43148),
            .I(N__43145));
    Span4Mux_v I__9555 (
            .O(N__43145),
            .I(N__43142));
    Odrv4 I__9554 (
            .O(N__43142),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt22 ));
    InMux I__9553 (
            .O(N__43139),
            .I(N__43136));
    LocalMux I__9552 (
            .O(N__43136),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    CascadeMux I__9551 (
            .O(N__43133),
            .I(N__43130));
    InMux I__9550 (
            .O(N__43130),
            .I(N__43127));
    LocalMux I__9549 (
            .O(N__43127),
            .I(N__43123));
    InMux I__9548 (
            .O(N__43126),
            .I(N__43120));
    Odrv4 I__9547 (
            .O(N__43123),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    LocalMux I__9546 (
            .O(N__43120),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    InMux I__9545 (
            .O(N__43115),
            .I(N__43112));
    LocalMux I__9544 (
            .O(N__43112),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__9543 (
            .O(N__43109),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ));
    InMux I__9542 (
            .O(N__43106),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    InMux I__9541 (
            .O(N__43103),
            .I(N__43099));
    InMux I__9540 (
            .O(N__43102),
            .I(N__43096));
    LocalMux I__9539 (
            .O(N__43099),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    LocalMux I__9538 (
            .O(N__43096),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    CascadeMux I__9537 (
            .O(N__43091),
            .I(N__43087));
    InMux I__9536 (
            .O(N__43090),
            .I(N__43084));
    InMux I__9535 (
            .O(N__43087),
            .I(N__43080));
    LocalMux I__9534 (
            .O(N__43084),
            .I(N__43077));
    InMux I__9533 (
            .O(N__43083),
            .I(N__43074));
    LocalMux I__9532 (
            .O(N__43080),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__9531 (
            .O(N__43077),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__9530 (
            .O(N__43074),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__9529 (
            .O(N__43067),
            .I(N__43064));
    InMux I__9528 (
            .O(N__43064),
            .I(N__43061));
    LocalMux I__9527 (
            .O(N__43061),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    InMux I__9526 (
            .O(N__43058),
            .I(N__43054));
    InMux I__9525 (
            .O(N__43057),
            .I(N__43051));
    LocalMux I__9524 (
            .O(N__43054),
            .I(N__43048));
    LocalMux I__9523 (
            .O(N__43051),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__9522 (
            .O(N__43048),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__9521 (
            .O(N__43043),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__9520 (
            .O(N__43040),
            .I(N__43037));
    LocalMux I__9519 (
            .O(N__43037),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ));
    CascadeMux I__9518 (
            .O(N__43034),
            .I(N__43030));
    InMux I__9517 (
            .O(N__43033),
            .I(N__43027));
    InMux I__9516 (
            .O(N__43030),
            .I(N__43024));
    LocalMux I__9515 (
            .O(N__43027),
            .I(N__43021));
    LocalMux I__9514 (
            .O(N__43024),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__9513 (
            .O(N__43021),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__9512 (
            .O(N__43016),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__9511 (
            .O(N__43013),
            .I(N__43010));
    LocalMux I__9510 (
            .O(N__43010),
            .I(N__43007));
    Span4Mux_v I__9509 (
            .O(N__43007),
            .I(N__43004));
    Odrv4 I__9508 (
            .O(N__43004),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__9507 (
            .O(N__43001),
            .I(N__42998));
    InMux I__9506 (
            .O(N__42998),
            .I(N__42995));
    LocalMux I__9505 (
            .O(N__42995),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__9504 (
            .O(N__42992),
            .I(N__42989));
    LocalMux I__9503 (
            .O(N__42989),
            .I(N__42986));
    Span4Mux_v I__9502 (
            .O(N__42986),
            .I(N__42983));
    Odrv4 I__9501 (
            .O(N__42983),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__9500 (
            .O(N__42980),
            .I(N__42977));
    InMux I__9499 (
            .O(N__42977),
            .I(N__42974));
    LocalMux I__9498 (
            .O(N__42974),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__9497 (
            .O(N__42971),
            .I(N__42968));
    InMux I__9496 (
            .O(N__42968),
            .I(N__42965));
    LocalMux I__9495 (
            .O(N__42965),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__9494 (
            .O(N__42962),
            .I(N__42959));
    InMux I__9493 (
            .O(N__42959),
            .I(N__42956));
    LocalMux I__9492 (
            .O(N__42956),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__9491 (
            .O(N__42953),
            .I(N__42950));
    LocalMux I__9490 (
            .O(N__42950),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__9489 (
            .O(N__42947),
            .I(N__42944));
    LocalMux I__9488 (
            .O(N__42944),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__9487 (
            .O(N__42941),
            .I(N__42938));
    InMux I__9486 (
            .O(N__42938),
            .I(N__42935));
    LocalMux I__9485 (
            .O(N__42935),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__9484 (
            .O(N__42932),
            .I(N__42929));
    LocalMux I__9483 (
            .O(N__42929),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__9482 (
            .O(N__42926),
            .I(N__42923));
    InMux I__9481 (
            .O(N__42923),
            .I(N__42920));
    LocalMux I__9480 (
            .O(N__42920),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__9479 (
            .O(N__42917),
            .I(N__42914));
    LocalMux I__9478 (
            .O(N__42914),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__9477 (
            .O(N__42911),
            .I(N__42908));
    InMux I__9476 (
            .O(N__42908),
            .I(N__42905));
    LocalMux I__9475 (
            .O(N__42905),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__9474 (
            .O(N__42902),
            .I(N__42899));
    LocalMux I__9473 (
            .O(N__42899),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__9472 (
            .O(N__42896),
            .I(N__42893));
    InMux I__9471 (
            .O(N__42893),
            .I(N__42890));
    LocalMux I__9470 (
            .O(N__42890),
            .I(N__42887));
    Odrv4 I__9469 (
            .O(N__42887),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__9468 (
            .O(N__42884),
            .I(N__42881));
    LocalMux I__9467 (
            .O(N__42881),
            .I(N__42878));
    Span4Mux_h I__9466 (
            .O(N__42878),
            .I(N__42875));
    Odrv4 I__9465 (
            .O(N__42875),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__9464 (
            .O(N__42872),
            .I(N__42869));
    InMux I__9463 (
            .O(N__42869),
            .I(N__42866));
    LocalMux I__9462 (
            .O(N__42866),
            .I(N__42863));
    Odrv4 I__9461 (
            .O(N__42863),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__9460 (
            .O(N__42860),
            .I(N__42857));
    LocalMux I__9459 (
            .O(N__42857),
            .I(N__42854));
    Span4Mux_h I__9458 (
            .O(N__42854),
            .I(N__42851));
    Odrv4 I__9457 (
            .O(N__42851),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__9456 (
            .O(N__42848),
            .I(N__42845));
    InMux I__9455 (
            .O(N__42845),
            .I(N__42842));
    LocalMux I__9454 (
            .O(N__42842),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__9453 (
            .O(N__42839),
            .I(N__42836));
    LocalMux I__9452 (
            .O(N__42836),
            .I(N__42833));
    Span4Mux_h I__9451 (
            .O(N__42833),
            .I(N__42830));
    Odrv4 I__9450 (
            .O(N__42830),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__9449 (
            .O(N__42827),
            .I(N__42824));
    InMux I__9448 (
            .O(N__42824),
            .I(N__42821));
    LocalMux I__9447 (
            .O(N__42821),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__9446 (
            .O(N__42818),
            .I(N__42815));
    LocalMux I__9445 (
            .O(N__42815),
            .I(N__42812));
    Odrv4 I__9444 (
            .O(N__42812),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__9443 (
            .O(N__42809),
            .I(N__42806));
    LocalMux I__9442 (
            .O(N__42806),
            .I(N__42803));
    Odrv4 I__9441 (
            .O(N__42803),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__9440 (
            .O(N__42800),
            .I(N__42797));
    LocalMux I__9439 (
            .O(N__42797),
            .I(N__42794));
    Odrv4 I__9438 (
            .O(N__42794),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    CascadeMux I__9437 (
            .O(N__42791),
            .I(N__42788));
    InMux I__9436 (
            .O(N__42788),
            .I(N__42785));
    LocalMux I__9435 (
            .O(N__42785),
            .I(N__42782));
    Odrv4 I__9434 (
            .O(N__42782),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__9433 (
            .O(N__42779),
            .I(N__42776));
    LocalMux I__9432 (
            .O(N__42776),
            .I(N__42773));
    Span4Mux_h I__9431 (
            .O(N__42773),
            .I(N__42770));
    Odrv4 I__9430 (
            .O(N__42770),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__9429 (
            .O(N__42767),
            .I(N__42764));
    LocalMux I__9428 (
            .O(N__42764),
            .I(N__42761));
    Odrv4 I__9427 (
            .O(N__42761),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__9426 (
            .O(N__42758),
            .I(N__42754));
    InMux I__9425 (
            .O(N__42757),
            .I(N__42750));
    LocalMux I__9424 (
            .O(N__42754),
            .I(N__42746));
    InMux I__9423 (
            .O(N__42753),
            .I(N__42743));
    LocalMux I__9422 (
            .O(N__42750),
            .I(N__42740));
    InMux I__9421 (
            .O(N__42749),
            .I(N__42737));
    Span4Mux_v I__9420 (
            .O(N__42746),
            .I(N__42734));
    LocalMux I__9419 (
            .O(N__42743),
            .I(N__42731));
    Span4Mux_v I__9418 (
            .O(N__42740),
            .I(N__42726));
    LocalMux I__9417 (
            .O(N__42737),
            .I(N__42726));
    Span4Mux_h I__9416 (
            .O(N__42734),
            .I(N__42723));
    Span4Mux_v I__9415 (
            .O(N__42731),
            .I(N__42720));
    Span4Mux_h I__9414 (
            .O(N__42726),
            .I(N__42715));
    Span4Mux_h I__9413 (
            .O(N__42723),
            .I(N__42715));
    Odrv4 I__9412 (
            .O(N__42720),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__9411 (
            .O(N__42715),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__9410 (
            .O(N__42710),
            .I(N__42707));
    InMux I__9409 (
            .O(N__42707),
            .I(N__42704));
    LocalMux I__9408 (
            .O(N__42704),
            .I(N__42701));
    Span4Mux_v I__9407 (
            .O(N__42701),
            .I(N__42698));
    Span4Mux_h I__9406 (
            .O(N__42698),
            .I(N__42695));
    Span4Mux_h I__9405 (
            .O(N__42695),
            .I(N__42692));
    Odrv4 I__9404 (
            .O(N__42692),
            .I(\current_shift_inst.PI_CTRL.integrator_i_29 ));
    CascadeMux I__9403 (
            .O(N__42689),
            .I(N__42686));
    InMux I__9402 (
            .O(N__42686),
            .I(N__42683));
    LocalMux I__9401 (
            .O(N__42683),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__9400 (
            .O(N__42680),
            .I(N__42677));
    InMux I__9399 (
            .O(N__42677),
            .I(N__42674));
    LocalMux I__9398 (
            .O(N__42674),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__9397 (
            .O(N__42671),
            .I(N__42668));
    LocalMux I__9396 (
            .O(N__42668),
            .I(N__42665));
    Odrv4 I__9395 (
            .O(N__42665),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    CascadeMux I__9394 (
            .O(N__42662),
            .I(N__42659));
    InMux I__9393 (
            .O(N__42659),
            .I(N__42656));
    LocalMux I__9392 (
            .O(N__42656),
            .I(N__42653));
    Odrv4 I__9391 (
            .O(N__42653),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__9390 (
            .O(N__42650),
            .I(N__42647));
    LocalMux I__9389 (
            .O(N__42647),
            .I(N__42644));
    Odrv4 I__9388 (
            .O(N__42644),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__9387 (
            .O(N__42641),
            .I(N__42638));
    LocalMux I__9386 (
            .O(N__42638),
            .I(N__42635));
    Odrv4 I__9385 (
            .O(N__42635),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    CascadeMux I__9384 (
            .O(N__42632),
            .I(N__42629));
    InMux I__9383 (
            .O(N__42629),
            .I(N__42626));
    LocalMux I__9382 (
            .O(N__42626),
            .I(N__42623));
    Odrv4 I__9381 (
            .O(N__42623),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__9380 (
            .O(N__42620),
            .I(N__42617));
    LocalMux I__9379 (
            .O(N__42617),
            .I(N__42614));
    Span4Mux_v I__9378 (
            .O(N__42614),
            .I(N__42611));
    Odrv4 I__9377 (
            .O(N__42611),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    CascadeMux I__9376 (
            .O(N__42608),
            .I(N__42605));
    InMux I__9375 (
            .O(N__42605),
            .I(N__42602));
    LocalMux I__9374 (
            .O(N__42602),
            .I(N__42599));
    Odrv4 I__9373 (
            .O(N__42599),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__9372 (
            .O(N__42596),
            .I(N__42593));
    LocalMux I__9371 (
            .O(N__42593),
            .I(N__42590));
    Span4Mux_h I__9370 (
            .O(N__42590),
            .I(N__42587));
    Odrv4 I__9369 (
            .O(N__42587),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__9368 (
            .O(N__42584),
            .I(N__42581));
    LocalMux I__9367 (
            .O(N__42581),
            .I(N__42578));
    Odrv4 I__9366 (
            .O(N__42578),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__9365 (
            .O(N__42575),
            .I(N__42572));
    LocalMux I__9364 (
            .O(N__42572),
            .I(N__42567));
    InMux I__9363 (
            .O(N__42571),
            .I(N__42564));
    InMux I__9362 (
            .O(N__42570),
            .I(N__42561));
    Span4Mux_v I__9361 (
            .O(N__42567),
            .I(N__42556));
    LocalMux I__9360 (
            .O(N__42564),
            .I(N__42556));
    LocalMux I__9359 (
            .O(N__42561),
            .I(N__42553));
    Odrv4 I__9358 (
            .O(N__42556),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__9357 (
            .O(N__42553),
            .I(\current_shift_inst.un4_control_input1_17 ));
    InMux I__9356 (
            .O(N__42548),
            .I(N__42543));
    InMux I__9355 (
            .O(N__42547),
            .I(N__42540));
    InMux I__9354 (
            .O(N__42546),
            .I(N__42537));
    LocalMux I__9353 (
            .O(N__42543),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__9352 (
            .O(N__42540),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__9351 (
            .O(N__42537),
            .I(\current_shift_inst.un4_control_input1_20 ));
    CascadeMux I__9350 (
            .O(N__42530),
            .I(N__42527));
    InMux I__9349 (
            .O(N__42527),
            .I(N__42524));
    LocalMux I__9348 (
            .O(N__42524),
            .I(N__42521));
    Span4Mux_h I__9347 (
            .O(N__42521),
            .I(N__42518));
    Odrv4 I__9346 (
            .O(N__42518),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    CascadeMux I__9345 (
            .O(N__42515),
            .I(N__42511));
    InMux I__9344 (
            .O(N__42514),
            .I(N__42507));
    InMux I__9343 (
            .O(N__42511),
            .I(N__42502));
    InMux I__9342 (
            .O(N__42510),
            .I(N__42502));
    LocalMux I__9341 (
            .O(N__42507),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__9340 (
            .O(N__42502),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__9339 (
            .O(N__42497),
            .I(N__42494));
    LocalMux I__9338 (
            .O(N__42494),
            .I(N__42491));
    Span4Mux_h I__9337 (
            .O(N__42491),
            .I(N__42488));
    Odrv4 I__9336 (
            .O(N__42488),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__9335 (
            .O(N__42485),
            .I(N__42482));
    LocalMux I__9334 (
            .O(N__42482),
            .I(N__42479));
    Odrv4 I__9333 (
            .O(N__42479),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    CascadeMux I__9332 (
            .O(N__42476),
            .I(N__42462));
    CascadeMux I__9331 (
            .O(N__42475),
            .I(N__42456));
    CascadeMux I__9330 (
            .O(N__42474),
            .I(N__42453));
    CascadeMux I__9329 (
            .O(N__42473),
            .I(N__42448));
    CascadeMux I__9328 (
            .O(N__42472),
            .I(N__42434));
    CascadeMux I__9327 (
            .O(N__42471),
            .I(N__42428));
    CascadeMux I__9326 (
            .O(N__42470),
            .I(N__42425));
    CascadeMux I__9325 (
            .O(N__42469),
            .I(N__42417));
    CascadeMux I__9324 (
            .O(N__42468),
            .I(N__42413));
    CascadeMux I__9323 (
            .O(N__42467),
            .I(N__42408));
    CascadeMux I__9322 (
            .O(N__42466),
            .I(N__42404));
    CascadeMux I__9321 (
            .O(N__42465),
            .I(N__42400));
    InMux I__9320 (
            .O(N__42462),
            .I(N__42384));
    InMux I__9319 (
            .O(N__42461),
            .I(N__42373));
    InMux I__9318 (
            .O(N__42460),
            .I(N__42373));
    InMux I__9317 (
            .O(N__42459),
            .I(N__42373));
    InMux I__9316 (
            .O(N__42456),
            .I(N__42373));
    InMux I__9315 (
            .O(N__42453),
            .I(N__42373));
    InMux I__9314 (
            .O(N__42452),
            .I(N__42370));
    InMux I__9313 (
            .O(N__42451),
            .I(N__42359));
    InMux I__9312 (
            .O(N__42448),
            .I(N__42359));
    InMux I__9311 (
            .O(N__42447),
            .I(N__42359));
    InMux I__9310 (
            .O(N__42446),
            .I(N__42359));
    InMux I__9309 (
            .O(N__42445),
            .I(N__42359));
    InMux I__9308 (
            .O(N__42444),
            .I(N__42342));
    InMux I__9307 (
            .O(N__42443),
            .I(N__42342));
    InMux I__9306 (
            .O(N__42442),
            .I(N__42342));
    InMux I__9305 (
            .O(N__42441),
            .I(N__42342));
    InMux I__9304 (
            .O(N__42440),
            .I(N__42342));
    InMux I__9303 (
            .O(N__42439),
            .I(N__42342));
    InMux I__9302 (
            .O(N__42438),
            .I(N__42342));
    InMux I__9301 (
            .O(N__42437),
            .I(N__42342));
    InMux I__9300 (
            .O(N__42434),
            .I(N__42339));
    InMux I__9299 (
            .O(N__42433),
            .I(N__42328));
    InMux I__9298 (
            .O(N__42432),
            .I(N__42328));
    InMux I__9297 (
            .O(N__42431),
            .I(N__42328));
    InMux I__9296 (
            .O(N__42428),
            .I(N__42328));
    InMux I__9295 (
            .O(N__42425),
            .I(N__42328));
    CascadeMux I__9294 (
            .O(N__42424),
            .I(N__42315));
    CascadeMux I__9293 (
            .O(N__42423),
            .I(N__42311));
    CascadeMux I__9292 (
            .O(N__42422),
            .I(N__42307));
    InMux I__9291 (
            .O(N__42421),
            .I(N__42291));
    InMux I__9290 (
            .O(N__42420),
            .I(N__42291));
    InMux I__9289 (
            .O(N__42417),
            .I(N__42274));
    InMux I__9288 (
            .O(N__42416),
            .I(N__42274));
    InMux I__9287 (
            .O(N__42413),
            .I(N__42274));
    InMux I__9286 (
            .O(N__42412),
            .I(N__42274));
    InMux I__9285 (
            .O(N__42411),
            .I(N__42274));
    InMux I__9284 (
            .O(N__42408),
            .I(N__42274));
    InMux I__9283 (
            .O(N__42407),
            .I(N__42274));
    InMux I__9282 (
            .O(N__42404),
            .I(N__42274));
    InMux I__9281 (
            .O(N__42403),
            .I(N__42265));
    InMux I__9280 (
            .O(N__42400),
            .I(N__42265));
    InMux I__9279 (
            .O(N__42399),
            .I(N__42265));
    InMux I__9278 (
            .O(N__42398),
            .I(N__42265));
    CascadeMux I__9277 (
            .O(N__42397),
            .I(N__42262));
    CascadeMux I__9276 (
            .O(N__42396),
            .I(N__42258));
    CascadeMux I__9275 (
            .O(N__42395),
            .I(N__42254));
    CascadeMux I__9274 (
            .O(N__42394),
            .I(N__42250));
    CascadeMux I__9273 (
            .O(N__42393),
            .I(N__42238));
    CascadeMux I__9272 (
            .O(N__42392),
            .I(N__42234));
    CascadeMux I__9271 (
            .O(N__42391),
            .I(N__42230));
    CascadeMux I__9270 (
            .O(N__42390),
            .I(N__42226));
    CascadeMux I__9269 (
            .O(N__42389),
            .I(N__42222));
    CascadeMux I__9268 (
            .O(N__42388),
            .I(N__42218));
    CascadeMux I__9267 (
            .O(N__42387),
            .I(N__42214));
    LocalMux I__9266 (
            .O(N__42384),
            .I(N__42208));
    LocalMux I__9265 (
            .O(N__42373),
            .I(N__42208));
    LocalMux I__9264 (
            .O(N__42370),
            .I(N__42205));
    LocalMux I__9263 (
            .O(N__42359),
            .I(N__42200));
    LocalMux I__9262 (
            .O(N__42342),
            .I(N__42200));
    LocalMux I__9261 (
            .O(N__42339),
            .I(N__42195));
    LocalMux I__9260 (
            .O(N__42328),
            .I(N__42195));
    InMux I__9259 (
            .O(N__42327),
            .I(N__42188));
    InMux I__9258 (
            .O(N__42326),
            .I(N__42188));
    InMux I__9257 (
            .O(N__42325),
            .I(N__42188));
    CascadeMux I__9256 (
            .O(N__42324),
            .I(N__42185));
    CascadeMux I__9255 (
            .O(N__42323),
            .I(N__42179));
    CascadeMux I__9254 (
            .O(N__42322),
            .I(N__42176));
    CascadeMux I__9253 (
            .O(N__42321),
            .I(N__42173));
    CascadeMux I__9252 (
            .O(N__42320),
            .I(N__42170));
    CascadeMux I__9251 (
            .O(N__42319),
            .I(N__42167));
    InMux I__9250 (
            .O(N__42318),
            .I(N__42145));
    InMux I__9249 (
            .O(N__42315),
            .I(N__42145));
    InMux I__9248 (
            .O(N__42314),
            .I(N__42145));
    InMux I__9247 (
            .O(N__42311),
            .I(N__42145));
    InMux I__9246 (
            .O(N__42310),
            .I(N__42145));
    InMux I__9245 (
            .O(N__42307),
            .I(N__42145));
    InMux I__9244 (
            .O(N__42306),
            .I(N__42145));
    CascadeMux I__9243 (
            .O(N__42305),
            .I(N__42140));
    CascadeMux I__9242 (
            .O(N__42304),
            .I(N__42136));
    CascadeMux I__9241 (
            .O(N__42303),
            .I(N__42132));
    CascadeMux I__9240 (
            .O(N__42302),
            .I(N__42128));
    CascadeMux I__9239 (
            .O(N__42301),
            .I(N__42124));
    CascadeMux I__9238 (
            .O(N__42300),
            .I(N__42120));
    CascadeMux I__9237 (
            .O(N__42299),
            .I(N__42116));
    CascadeMux I__9236 (
            .O(N__42298),
            .I(N__42112));
    CascadeMux I__9235 (
            .O(N__42297),
            .I(N__42108));
    CascadeMux I__9234 (
            .O(N__42296),
            .I(N__42104));
    LocalMux I__9233 (
            .O(N__42291),
            .I(N__42096));
    LocalMux I__9232 (
            .O(N__42274),
            .I(N__42096));
    LocalMux I__9231 (
            .O(N__42265),
            .I(N__42096));
    InMux I__9230 (
            .O(N__42262),
            .I(N__42079));
    InMux I__9229 (
            .O(N__42261),
            .I(N__42079));
    InMux I__9228 (
            .O(N__42258),
            .I(N__42079));
    InMux I__9227 (
            .O(N__42257),
            .I(N__42079));
    InMux I__9226 (
            .O(N__42254),
            .I(N__42079));
    InMux I__9225 (
            .O(N__42253),
            .I(N__42079));
    InMux I__9224 (
            .O(N__42250),
            .I(N__42079));
    InMux I__9223 (
            .O(N__42249),
            .I(N__42079));
    InMux I__9222 (
            .O(N__42248),
            .I(N__42070));
    InMux I__9221 (
            .O(N__42247),
            .I(N__42070));
    InMux I__9220 (
            .O(N__42246),
            .I(N__42070));
    InMux I__9219 (
            .O(N__42245),
            .I(N__42070));
    InMux I__9218 (
            .O(N__42244),
            .I(N__42061));
    InMux I__9217 (
            .O(N__42243),
            .I(N__42061));
    InMux I__9216 (
            .O(N__42242),
            .I(N__42061));
    InMux I__9215 (
            .O(N__42241),
            .I(N__42061));
    InMux I__9214 (
            .O(N__42238),
            .I(N__42044));
    InMux I__9213 (
            .O(N__42237),
            .I(N__42044));
    InMux I__9212 (
            .O(N__42234),
            .I(N__42044));
    InMux I__9211 (
            .O(N__42233),
            .I(N__42044));
    InMux I__9210 (
            .O(N__42230),
            .I(N__42044));
    InMux I__9209 (
            .O(N__42229),
            .I(N__42044));
    InMux I__9208 (
            .O(N__42226),
            .I(N__42044));
    InMux I__9207 (
            .O(N__42225),
            .I(N__42044));
    InMux I__9206 (
            .O(N__42222),
            .I(N__42031));
    InMux I__9205 (
            .O(N__42221),
            .I(N__42031));
    InMux I__9204 (
            .O(N__42218),
            .I(N__42031));
    InMux I__9203 (
            .O(N__42217),
            .I(N__42031));
    InMux I__9202 (
            .O(N__42214),
            .I(N__42031));
    InMux I__9201 (
            .O(N__42213),
            .I(N__42031));
    Span12Mux_s11_h I__9200 (
            .O(N__42208),
            .I(N__42028));
    Span4Mux_v I__9199 (
            .O(N__42205),
            .I(N__42019));
    Span4Mux_h I__9198 (
            .O(N__42200),
            .I(N__42019));
    Span4Mux_v I__9197 (
            .O(N__42195),
            .I(N__42019));
    LocalMux I__9196 (
            .O(N__42188),
            .I(N__42019));
    InMux I__9195 (
            .O(N__42185),
            .I(N__42010));
    InMux I__9194 (
            .O(N__42184),
            .I(N__42010));
    InMux I__9193 (
            .O(N__42183),
            .I(N__42010));
    InMux I__9192 (
            .O(N__42182),
            .I(N__42010));
    InMux I__9191 (
            .O(N__42179),
            .I(N__42003));
    InMux I__9190 (
            .O(N__42176),
            .I(N__42003));
    InMux I__9189 (
            .O(N__42173),
            .I(N__42003));
    InMux I__9188 (
            .O(N__42170),
            .I(N__42000));
    InMux I__9187 (
            .O(N__42167),
            .I(N__41985));
    InMux I__9186 (
            .O(N__42166),
            .I(N__41985));
    InMux I__9185 (
            .O(N__42165),
            .I(N__41985));
    InMux I__9184 (
            .O(N__42164),
            .I(N__41985));
    InMux I__9183 (
            .O(N__42163),
            .I(N__41985));
    InMux I__9182 (
            .O(N__42162),
            .I(N__41985));
    InMux I__9181 (
            .O(N__42161),
            .I(N__41985));
    InMux I__9180 (
            .O(N__42160),
            .I(N__41982));
    LocalMux I__9179 (
            .O(N__42145),
            .I(N__41979));
    InMux I__9178 (
            .O(N__42144),
            .I(N__41962));
    InMux I__9177 (
            .O(N__42143),
            .I(N__41962));
    InMux I__9176 (
            .O(N__42140),
            .I(N__41962));
    InMux I__9175 (
            .O(N__42139),
            .I(N__41962));
    InMux I__9174 (
            .O(N__42136),
            .I(N__41962));
    InMux I__9173 (
            .O(N__42135),
            .I(N__41962));
    InMux I__9172 (
            .O(N__42132),
            .I(N__41962));
    InMux I__9171 (
            .O(N__42131),
            .I(N__41962));
    InMux I__9170 (
            .O(N__42128),
            .I(N__41945));
    InMux I__9169 (
            .O(N__42127),
            .I(N__41945));
    InMux I__9168 (
            .O(N__42124),
            .I(N__41945));
    InMux I__9167 (
            .O(N__42123),
            .I(N__41945));
    InMux I__9166 (
            .O(N__42120),
            .I(N__41945));
    InMux I__9165 (
            .O(N__42119),
            .I(N__41945));
    InMux I__9164 (
            .O(N__42116),
            .I(N__41945));
    InMux I__9163 (
            .O(N__42115),
            .I(N__41945));
    InMux I__9162 (
            .O(N__42112),
            .I(N__41932));
    InMux I__9161 (
            .O(N__42111),
            .I(N__41932));
    InMux I__9160 (
            .O(N__42108),
            .I(N__41932));
    InMux I__9159 (
            .O(N__42107),
            .I(N__41932));
    InMux I__9158 (
            .O(N__42104),
            .I(N__41932));
    InMux I__9157 (
            .O(N__42103),
            .I(N__41932));
    Span12Mux_s11_h I__9156 (
            .O(N__42096),
            .I(N__41919));
    LocalMux I__9155 (
            .O(N__42079),
            .I(N__41919));
    LocalMux I__9154 (
            .O(N__42070),
            .I(N__41919));
    LocalMux I__9153 (
            .O(N__42061),
            .I(N__41919));
    LocalMux I__9152 (
            .O(N__42044),
            .I(N__41919));
    LocalMux I__9151 (
            .O(N__42031),
            .I(N__41919));
    Odrv12 I__9150 (
            .O(N__42028),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__9149 (
            .O(N__42019),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9148 (
            .O(N__42010),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9147 (
            .O(N__42003),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9146 (
            .O(N__42000),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9145 (
            .O(N__41985),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9144 (
            .O(N__41982),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__9143 (
            .O(N__41979),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9142 (
            .O(N__41962),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9141 (
            .O(N__41945),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9140 (
            .O(N__41932),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__9139 (
            .O(N__41919),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__9138 (
            .O(N__41894),
            .I(N__41891));
    InMux I__9137 (
            .O(N__41891),
            .I(N__41888));
    LocalMux I__9136 (
            .O(N__41888),
            .I(N__41885));
    Span4Mux_h I__9135 (
            .O(N__41885),
            .I(N__41882));
    Odrv4 I__9134 (
            .O(N__41882),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    CascadeMux I__9133 (
            .O(N__41879),
            .I(N__41875));
    InMux I__9132 (
            .O(N__41878),
            .I(N__41867));
    InMux I__9131 (
            .O(N__41875),
            .I(N__41867));
    InMux I__9130 (
            .O(N__41874),
            .I(N__41867));
    LocalMux I__9129 (
            .O(N__41867),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__9128 (
            .O(N__41864),
            .I(N__41849));
    InMux I__9127 (
            .O(N__41863),
            .I(N__41840));
    InMux I__9126 (
            .O(N__41862),
            .I(N__41827));
    InMux I__9125 (
            .O(N__41861),
            .I(N__41827));
    InMux I__9124 (
            .O(N__41860),
            .I(N__41827));
    InMux I__9123 (
            .O(N__41859),
            .I(N__41827));
    InMux I__9122 (
            .O(N__41858),
            .I(N__41827));
    InMux I__9121 (
            .O(N__41857),
            .I(N__41827));
    InMux I__9120 (
            .O(N__41856),
            .I(N__41816));
    InMux I__9119 (
            .O(N__41855),
            .I(N__41816));
    InMux I__9118 (
            .O(N__41854),
            .I(N__41816));
    InMux I__9117 (
            .O(N__41853),
            .I(N__41816));
    InMux I__9116 (
            .O(N__41852),
            .I(N__41816));
    LocalMux I__9115 (
            .O(N__41849),
            .I(N__41813));
    InMux I__9114 (
            .O(N__41848),
            .I(N__41808));
    InMux I__9113 (
            .O(N__41847),
            .I(N__41808));
    InMux I__9112 (
            .O(N__41846),
            .I(N__41793));
    InMux I__9111 (
            .O(N__41845),
            .I(N__41793));
    InMux I__9110 (
            .O(N__41844),
            .I(N__41793));
    InMux I__9109 (
            .O(N__41843),
            .I(N__41793));
    LocalMux I__9108 (
            .O(N__41840),
            .I(N__41786));
    LocalMux I__9107 (
            .O(N__41827),
            .I(N__41786));
    LocalMux I__9106 (
            .O(N__41816),
            .I(N__41786));
    Span4Mux_v I__9105 (
            .O(N__41813),
            .I(N__41781));
    LocalMux I__9104 (
            .O(N__41808),
            .I(N__41781));
    InMux I__9103 (
            .O(N__41807),
            .I(N__41778));
    InMux I__9102 (
            .O(N__41806),
            .I(N__41767));
    InMux I__9101 (
            .O(N__41805),
            .I(N__41767));
    InMux I__9100 (
            .O(N__41804),
            .I(N__41767));
    InMux I__9099 (
            .O(N__41803),
            .I(N__41767));
    InMux I__9098 (
            .O(N__41802),
            .I(N__41767));
    LocalMux I__9097 (
            .O(N__41793),
            .I(N__41760));
    Span4Mux_v I__9096 (
            .O(N__41786),
            .I(N__41760));
    Span4Mux_h I__9095 (
            .O(N__41781),
            .I(N__41760));
    LocalMux I__9094 (
            .O(N__41778),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__9093 (
            .O(N__41767),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__9092 (
            .O(N__41760),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__9091 (
            .O(N__41753),
            .I(N__41750));
    LocalMux I__9090 (
            .O(N__41750),
            .I(N__41745));
    InMux I__9089 (
            .O(N__41749),
            .I(N__41742));
    InMux I__9088 (
            .O(N__41748),
            .I(N__41739));
    Odrv4 I__9087 (
            .O(N__41745),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__9086 (
            .O(N__41742),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__9085 (
            .O(N__41739),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__9084 (
            .O(N__41732),
            .I(N__41729));
    LocalMux I__9083 (
            .O(N__41729),
            .I(N__41724));
    InMux I__9082 (
            .O(N__41728),
            .I(N__41721));
    InMux I__9081 (
            .O(N__41727),
            .I(N__41718));
    Odrv4 I__9080 (
            .O(N__41724),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__9079 (
            .O(N__41721),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__9078 (
            .O(N__41718),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__9077 (
            .O(N__41711),
            .I(N__41708));
    LocalMux I__9076 (
            .O(N__41708),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    CascadeMux I__9075 (
            .O(N__41705),
            .I(N__41702));
    InMux I__9074 (
            .O(N__41702),
            .I(N__41699));
    LocalMux I__9073 (
            .O(N__41699),
            .I(N__41695));
    InMux I__9072 (
            .O(N__41698),
            .I(N__41691));
    Span4Mux_h I__9071 (
            .O(N__41695),
            .I(N__41688));
    InMux I__9070 (
            .O(N__41694),
            .I(N__41685));
    LocalMux I__9069 (
            .O(N__41691),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__9068 (
            .O(N__41688),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__9067 (
            .O(N__41685),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__9066 (
            .O(N__41678),
            .I(N__41673));
    InMux I__9065 (
            .O(N__41677),
            .I(N__41670));
    InMux I__9064 (
            .O(N__41676),
            .I(N__41667));
    LocalMux I__9063 (
            .O(N__41673),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__9062 (
            .O(N__41670),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__9061 (
            .O(N__41667),
            .I(\current_shift_inst.un4_control_input1_18 ));
    CascadeMux I__9060 (
            .O(N__41660),
            .I(N__41657));
    InMux I__9059 (
            .O(N__41657),
            .I(N__41654));
    LocalMux I__9058 (
            .O(N__41654),
            .I(N__41650));
    InMux I__9057 (
            .O(N__41653),
            .I(N__41647));
    Span4Mux_v I__9056 (
            .O(N__41650),
            .I(N__41641));
    LocalMux I__9055 (
            .O(N__41647),
            .I(N__41641));
    InMux I__9054 (
            .O(N__41646),
            .I(N__41638));
    Odrv4 I__9053 (
            .O(N__41641),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__9052 (
            .O(N__41638),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__9051 (
            .O(N__41633),
            .I(N__41630));
    LocalMux I__9050 (
            .O(N__41630),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__9049 (
            .O(N__41627),
            .I(N__41624));
    LocalMux I__9048 (
            .O(N__41624),
            .I(N__41619));
    InMux I__9047 (
            .O(N__41623),
            .I(N__41616));
    InMux I__9046 (
            .O(N__41622),
            .I(N__41613));
    Odrv12 I__9045 (
            .O(N__41619),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__9044 (
            .O(N__41616),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__9043 (
            .O(N__41613),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__9042 (
            .O(N__41606),
            .I(N__41603));
    LocalMux I__9041 (
            .O(N__41603),
            .I(N__41599));
    InMux I__9040 (
            .O(N__41602),
            .I(N__41595));
    Span4Mux_h I__9039 (
            .O(N__41599),
            .I(N__41592));
    InMux I__9038 (
            .O(N__41598),
            .I(N__41589));
    LocalMux I__9037 (
            .O(N__41595),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__9036 (
            .O(N__41592),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__9035 (
            .O(N__41589),
            .I(\current_shift_inst.un4_control_input1_28 ));
    CascadeMux I__9034 (
            .O(N__41582),
            .I(N__41579));
    InMux I__9033 (
            .O(N__41579),
            .I(N__41576));
    LocalMux I__9032 (
            .O(N__41576),
            .I(N__41573));
    Span4Mux_v I__9031 (
            .O(N__41573),
            .I(N__41569));
    InMux I__9030 (
            .O(N__41572),
            .I(N__41566));
    Span4Mux_h I__9029 (
            .O(N__41569),
            .I(N__41562));
    LocalMux I__9028 (
            .O(N__41566),
            .I(N__41559));
    InMux I__9027 (
            .O(N__41565),
            .I(N__41556));
    Odrv4 I__9026 (
            .O(N__41562),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__9025 (
            .O(N__41559),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__9024 (
            .O(N__41556),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__9023 (
            .O(N__41549),
            .I(N__41546));
    LocalMux I__9022 (
            .O(N__41546),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    CascadeMux I__9021 (
            .O(N__41543),
            .I(N__41539));
    InMux I__9020 (
            .O(N__41542),
            .I(N__41536));
    InMux I__9019 (
            .O(N__41539),
            .I(N__41533));
    LocalMux I__9018 (
            .O(N__41536),
            .I(N__41529));
    LocalMux I__9017 (
            .O(N__41533),
            .I(N__41526));
    InMux I__9016 (
            .O(N__41532),
            .I(N__41523));
    Odrv4 I__9015 (
            .O(N__41529),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__9014 (
            .O(N__41526),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__9013 (
            .O(N__41523),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__9012 (
            .O(N__41516),
            .I(N__41512));
    InMux I__9011 (
            .O(N__41515),
            .I(N__41509));
    LocalMux I__9010 (
            .O(N__41512),
            .I(N__41503));
    LocalMux I__9009 (
            .O(N__41509),
            .I(N__41503));
    InMux I__9008 (
            .O(N__41508),
            .I(N__41500));
    Odrv4 I__9007 (
            .O(N__41503),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__9006 (
            .O(N__41500),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__9005 (
            .O(N__41495),
            .I(N__41492));
    LocalMux I__9004 (
            .O(N__41492),
            .I(N__41487));
    InMux I__9003 (
            .O(N__41491),
            .I(N__41484));
    InMux I__9002 (
            .O(N__41490),
            .I(N__41481));
    Odrv4 I__9001 (
            .O(N__41487),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__9000 (
            .O(N__41484),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__8999 (
            .O(N__41481),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__8998 (
            .O(N__41474),
            .I(N__41471));
    LocalMux I__8997 (
            .O(N__41471),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__8996 (
            .O(N__41468),
            .I(N__41464));
    InMux I__8995 (
            .O(N__41467),
            .I(N__41461));
    LocalMux I__8994 (
            .O(N__41464),
            .I(N__41457));
    LocalMux I__8993 (
            .O(N__41461),
            .I(N__41454));
    InMux I__8992 (
            .O(N__41460),
            .I(N__41451));
    Odrv4 I__8991 (
            .O(N__41457),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__8990 (
            .O(N__41454),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__8989 (
            .O(N__41451),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__8988 (
            .O(N__41444),
            .I(N__41441));
    LocalMux I__8987 (
            .O(N__41441),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__8986 (
            .O(N__41438),
            .I(N__41435));
    LocalMux I__8985 (
            .O(N__41435),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    CascadeMux I__8984 (
            .O(N__41432),
            .I(N__41429));
    InMux I__8983 (
            .O(N__41429),
            .I(N__41426));
    LocalMux I__8982 (
            .O(N__41426),
            .I(N__41421));
    InMux I__8981 (
            .O(N__41425),
            .I(N__41416));
    InMux I__8980 (
            .O(N__41424),
            .I(N__41416));
    Odrv4 I__8979 (
            .O(N__41421),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__8978 (
            .O(N__41416),
            .I(\current_shift_inst.un4_control_input1_8 ));
    CascadeMux I__8977 (
            .O(N__41411),
            .I(N__41408));
    InMux I__8976 (
            .O(N__41408),
            .I(N__41404));
    InMux I__8975 (
            .O(N__41407),
            .I(N__41401));
    LocalMux I__8974 (
            .O(N__41404),
            .I(N__41397));
    LocalMux I__8973 (
            .O(N__41401),
            .I(N__41394));
    InMux I__8972 (
            .O(N__41400),
            .I(N__41391));
    Odrv12 I__8971 (
            .O(N__41397),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__8970 (
            .O(N__41394),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__8969 (
            .O(N__41391),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__8968 (
            .O(N__41384),
            .I(N__41381));
    LocalMux I__8967 (
            .O(N__41381),
            .I(N__41376));
    InMux I__8966 (
            .O(N__41380),
            .I(N__41373));
    InMux I__8965 (
            .O(N__41379),
            .I(N__41370));
    Odrv4 I__8964 (
            .O(N__41376),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__8963 (
            .O(N__41373),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__8962 (
            .O(N__41370),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__8961 (
            .O(N__41363),
            .I(N__41359));
    InMux I__8960 (
            .O(N__41362),
            .I(N__41356));
    LocalMux I__8959 (
            .O(N__41359),
            .I(N__41353));
    LocalMux I__8958 (
            .O(N__41356),
            .I(N__41348));
    Span4Mux_h I__8957 (
            .O(N__41353),
            .I(N__41345));
    InMux I__8956 (
            .O(N__41352),
            .I(N__41340));
    InMux I__8955 (
            .O(N__41351),
            .I(N__41340));
    Odrv12 I__8954 (
            .O(N__41348),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    Odrv4 I__8953 (
            .O(N__41345),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__8952 (
            .O(N__41340),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__8951 (
            .O(N__41333),
            .I(N__41329));
    InMux I__8950 (
            .O(N__41332),
            .I(N__41326));
    LocalMux I__8949 (
            .O(N__41329),
            .I(N__41322));
    LocalMux I__8948 (
            .O(N__41326),
            .I(N__41319));
    InMux I__8947 (
            .O(N__41325),
            .I(N__41316));
    Odrv4 I__8946 (
            .O(N__41322),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__8945 (
            .O(N__41319),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__8944 (
            .O(N__41316),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__8943 (
            .O(N__41309),
            .I(N__41305));
    InMux I__8942 (
            .O(N__41308),
            .I(N__41302));
    LocalMux I__8941 (
            .O(N__41305),
            .I(N__41298));
    LocalMux I__8940 (
            .O(N__41302),
            .I(N__41295));
    InMux I__8939 (
            .O(N__41301),
            .I(N__41292));
    Odrv4 I__8938 (
            .O(N__41298),
            .I(\current_shift_inst.un4_control_input1_9 ));
    Odrv4 I__8937 (
            .O(N__41295),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__8936 (
            .O(N__41292),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__8935 (
            .O(N__41285),
            .I(N__41280));
    CascadeMux I__8934 (
            .O(N__41284),
            .I(N__41277));
    InMux I__8933 (
            .O(N__41283),
            .I(N__41273));
    LocalMux I__8932 (
            .O(N__41280),
            .I(N__41270));
    InMux I__8931 (
            .O(N__41277),
            .I(N__41267));
    InMux I__8930 (
            .O(N__41276),
            .I(N__41263));
    LocalMux I__8929 (
            .O(N__41273),
            .I(N__41260));
    Span4Mux_v I__8928 (
            .O(N__41270),
            .I(N__41257));
    LocalMux I__8927 (
            .O(N__41267),
            .I(N__41254));
    InMux I__8926 (
            .O(N__41266),
            .I(N__41251));
    LocalMux I__8925 (
            .O(N__41263),
            .I(N__41248));
    Span4Mux_v I__8924 (
            .O(N__41260),
            .I(N__41245));
    Span4Mux_h I__8923 (
            .O(N__41257),
            .I(N__41242));
    Span4Mux_h I__8922 (
            .O(N__41254),
            .I(N__41237));
    LocalMux I__8921 (
            .O(N__41251),
            .I(N__41237));
    Span4Mux_v I__8920 (
            .O(N__41248),
            .I(N__41230));
    Span4Mux_h I__8919 (
            .O(N__41245),
            .I(N__41230));
    Span4Mux_h I__8918 (
            .O(N__41242),
            .I(N__41230));
    Odrv4 I__8917 (
            .O(N__41237),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__8916 (
            .O(N__41230),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__8915 (
            .O(N__41225),
            .I(N__41222));
    LocalMux I__8914 (
            .O(N__41222),
            .I(N__41219));
    Span4Mux_v I__8913 (
            .O(N__41219),
            .I(N__41216));
    Sp12to4 I__8912 (
            .O(N__41216),
            .I(N__41213));
    Span12Mux_h I__8911 (
            .O(N__41213),
            .I(N__41210));
    Odrv12 I__8910 (
            .O(N__41210),
            .I(\current_shift_inst.PI_CTRL.integrator_i_11 ));
    CascadeMux I__8909 (
            .O(N__41207),
            .I(N__41204));
    InMux I__8908 (
            .O(N__41204),
            .I(N__41200));
    InMux I__8907 (
            .O(N__41203),
            .I(N__41196));
    LocalMux I__8906 (
            .O(N__41200),
            .I(N__41193));
    InMux I__8905 (
            .O(N__41199),
            .I(N__41190));
    LocalMux I__8904 (
            .O(N__41196),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__8903 (
            .O(N__41193),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__8902 (
            .O(N__41190),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__8901 (
            .O(N__41183),
            .I(N__41176));
    InMux I__8900 (
            .O(N__41182),
            .I(N__41176));
    InMux I__8899 (
            .O(N__41181),
            .I(N__41173));
    LocalMux I__8898 (
            .O(N__41176),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__8897 (
            .O(N__41173),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__8896 (
            .O(N__41168),
            .I(N__41164));
    InMux I__8895 (
            .O(N__41167),
            .I(N__41161));
    LocalMux I__8894 (
            .O(N__41164),
            .I(N__41157));
    LocalMux I__8893 (
            .O(N__41161),
            .I(N__41154));
    InMux I__8892 (
            .O(N__41160),
            .I(N__41151));
    Odrv4 I__8891 (
            .O(N__41157),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv12 I__8890 (
            .O(N__41154),
            .I(\current_shift_inst.un4_control_input1_16 ));
    LocalMux I__8889 (
            .O(N__41151),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__8888 (
            .O(N__41144),
            .I(N__41141));
    LocalMux I__8887 (
            .O(N__41141),
            .I(N__41137));
    InMux I__8886 (
            .O(N__41140),
            .I(N__41134));
    Span4Mux_h I__8885 (
            .O(N__41137),
            .I(N__41131));
    LocalMux I__8884 (
            .O(N__41134),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv4 I__8883 (
            .O(N__41131),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__8882 (
            .O(N__41126),
            .I(N__41123));
    InMux I__8881 (
            .O(N__41123),
            .I(N__41118));
    InMux I__8880 (
            .O(N__41122),
            .I(N__41115));
    InMux I__8879 (
            .O(N__41121),
            .I(N__41112));
    LocalMux I__8878 (
            .O(N__41118),
            .I(N__41107));
    LocalMux I__8877 (
            .O(N__41115),
            .I(N__41107));
    LocalMux I__8876 (
            .O(N__41112),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv4 I__8875 (
            .O(N__41107),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__8874 (
            .O(N__41102),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__8873 (
            .O(N__41099),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__8872 (
            .O(N__41096),
            .I(N__41091));
    CEMux I__8871 (
            .O(N__41095),
            .I(N__41088));
    CEMux I__8870 (
            .O(N__41094),
            .I(N__41084));
    LocalMux I__8869 (
            .O(N__41091),
            .I(N__41080));
    LocalMux I__8868 (
            .O(N__41088),
            .I(N__41077));
    CEMux I__8867 (
            .O(N__41087),
            .I(N__41074));
    LocalMux I__8866 (
            .O(N__41084),
            .I(N__41071));
    CEMux I__8865 (
            .O(N__41083),
            .I(N__41068));
    Span4Mux_v I__8864 (
            .O(N__41080),
            .I(N__41061));
    Span4Mux_v I__8863 (
            .O(N__41077),
            .I(N__41061));
    LocalMux I__8862 (
            .O(N__41074),
            .I(N__41061));
    Span4Mux_v I__8861 (
            .O(N__41071),
            .I(N__41058));
    LocalMux I__8860 (
            .O(N__41068),
            .I(N__41055));
    Span4Mux_v I__8859 (
            .O(N__41061),
            .I(N__41052));
    Span4Mux_v I__8858 (
            .O(N__41058),
            .I(N__41049));
    Span4Mux_v I__8857 (
            .O(N__41055),
            .I(N__41046));
    Span4Mux_h I__8856 (
            .O(N__41052),
            .I(N__41043));
    Odrv4 I__8855 (
            .O(N__41049),
            .I(\delay_measurement_inst.delay_hc_timer.N_201_i ));
    Odrv4 I__8854 (
            .O(N__41046),
            .I(\delay_measurement_inst.delay_hc_timer.N_201_i ));
    Odrv4 I__8853 (
            .O(N__41043),
            .I(\delay_measurement_inst.delay_hc_timer.N_201_i ));
    InMux I__8852 (
            .O(N__41036),
            .I(N__41030));
    InMux I__8851 (
            .O(N__41035),
            .I(N__41030));
    LocalMux I__8850 (
            .O(N__41030),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__8849 (
            .O(N__41027),
            .I(N__41024));
    LocalMux I__8848 (
            .O(N__41024),
            .I(N__41020));
    InMux I__8847 (
            .O(N__41023),
            .I(N__41017));
    Span4Mux_h I__8846 (
            .O(N__41020),
            .I(N__41011));
    LocalMux I__8845 (
            .O(N__41017),
            .I(N__41011));
    InMux I__8844 (
            .O(N__41016),
            .I(N__41008));
    Span4Mux_v I__8843 (
            .O(N__41011),
            .I(N__41002));
    LocalMux I__8842 (
            .O(N__41008),
            .I(N__41002));
    InMux I__8841 (
            .O(N__41007),
            .I(N__40999));
    Span4Mux_h I__8840 (
            .O(N__41002),
            .I(N__40996));
    LocalMux I__8839 (
            .O(N__40999),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__8838 (
            .O(N__40996),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__8837 (
            .O(N__40991),
            .I(N__40987));
    InMux I__8836 (
            .O(N__40990),
            .I(N__40983));
    LocalMux I__8835 (
            .O(N__40987),
            .I(N__40980));
    InMux I__8834 (
            .O(N__40986),
            .I(N__40977));
    LocalMux I__8833 (
            .O(N__40983),
            .I(N__40974));
    Span4Mux_v I__8832 (
            .O(N__40980),
            .I(N__40971));
    LocalMux I__8831 (
            .O(N__40977),
            .I(N__40966));
    Span4Mux_v I__8830 (
            .O(N__40974),
            .I(N__40966));
    Odrv4 I__8829 (
            .O(N__40971),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__8828 (
            .O(N__40966),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__8827 (
            .O(N__40961),
            .I(N__40956));
    InMux I__8826 (
            .O(N__40960),
            .I(N__40953));
    InMux I__8825 (
            .O(N__40959),
            .I(N__40950));
    LocalMux I__8824 (
            .O(N__40956),
            .I(N__40945));
    LocalMux I__8823 (
            .O(N__40953),
            .I(N__40945));
    LocalMux I__8822 (
            .O(N__40950),
            .I(N__40942));
    Span4Mux_v I__8821 (
            .O(N__40945),
            .I(N__40939));
    Span4Mux_v I__8820 (
            .O(N__40942),
            .I(N__40936));
    Odrv4 I__8819 (
            .O(N__40939),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    Odrv4 I__8818 (
            .O(N__40936),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    CascadeMux I__8817 (
            .O(N__40931),
            .I(N__40927));
    InMux I__8816 (
            .O(N__40930),
            .I(N__40922));
    InMux I__8815 (
            .O(N__40927),
            .I(N__40922));
    LocalMux I__8814 (
            .O(N__40922),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ));
    InMux I__8813 (
            .O(N__40919),
            .I(N__40916));
    LocalMux I__8812 (
            .O(N__40916),
            .I(N__40912));
    InMux I__8811 (
            .O(N__40915),
            .I(N__40909));
    Span4Mux_v I__8810 (
            .O(N__40912),
            .I(N__40905));
    LocalMux I__8809 (
            .O(N__40909),
            .I(N__40902));
    InMux I__8808 (
            .O(N__40908),
            .I(N__40899));
    Span4Mux_h I__8807 (
            .O(N__40905),
            .I(N__40894));
    Span4Mux_h I__8806 (
            .O(N__40902),
            .I(N__40894));
    LocalMux I__8805 (
            .O(N__40899),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    Odrv4 I__8804 (
            .O(N__40894),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    InMux I__8803 (
            .O(N__40889),
            .I(N__40884));
    InMux I__8802 (
            .O(N__40888),
            .I(N__40881));
    InMux I__8801 (
            .O(N__40887),
            .I(N__40878));
    LocalMux I__8800 (
            .O(N__40884),
            .I(N__40875));
    LocalMux I__8799 (
            .O(N__40881),
            .I(N__40868));
    LocalMux I__8798 (
            .O(N__40878),
            .I(N__40868));
    Span4Mux_h I__8797 (
            .O(N__40875),
            .I(N__40868));
    Odrv4 I__8796 (
            .O(N__40868),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    InMux I__8795 (
            .O(N__40865),
            .I(N__40859));
    InMux I__8794 (
            .O(N__40864),
            .I(N__40859));
    LocalMux I__8793 (
            .O(N__40859),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ));
    CascadeMux I__8792 (
            .O(N__40856),
            .I(N__40853));
    InMux I__8791 (
            .O(N__40853),
            .I(N__40850));
    LocalMux I__8790 (
            .O(N__40850),
            .I(N__40847));
    Odrv4 I__8789 (
            .O(N__40847),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    InMux I__8788 (
            .O(N__40844),
            .I(N__40841));
    LocalMux I__8787 (
            .O(N__40841),
            .I(N__40838));
    Span4Mux_h I__8786 (
            .O(N__40838),
            .I(N__40835));
    Odrv4 I__8785 (
            .O(N__40835),
            .I(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ));
    CascadeMux I__8784 (
            .O(N__40832),
            .I(N__40829));
    InMux I__8783 (
            .O(N__40829),
            .I(N__40824));
    InMux I__8782 (
            .O(N__40828),
            .I(N__40821));
    InMux I__8781 (
            .O(N__40827),
            .I(N__40818));
    LocalMux I__8780 (
            .O(N__40824),
            .I(N__40813));
    LocalMux I__8779 (
            .O(N__40821),
            .I(N__40813));
    LocalMux I__8778 (
            .O(N__40818),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv4 I__8777 (
            .O(N__40813),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__8776 (
            .O(N__40808),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__8775 (
            .O(N__40805),
            .I(N__40798));
    InMux I__8774 (
            .O(N__40804),
            .I(N__40798));
    InMux I__8773 (
            .O(N__40803),
            .I(N__40795));
    LocalMux I__8772 (
            .O(N__40798),
            .I(N__40792));
    LocalMux I__8771 (
            .O(N__40795),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv4 I__8770 (
            .O(N__40792),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__8769 (
            .O(N__40787),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__8768 (
            .O(N__40784),
            .I(N__40778));
    InMux I__8767 (
            .O(N__40783),
            .I(N__40778));
    LocalMux I__8766 (
            .O(N__40778),
            .I(N__40774));
    InMux I__8765 (
            .O(N__40777),
            .I(N__40771));
    Span4Mux_h I__8764 (
            .O(N__40774),
            .I(N__40768));
    LocalMux I__8763 (
            .O(N__40771),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv4 I__8762 (
            .O(N__40768),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__8761 (
            .O(N__40763),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__8760 (
            .O(N__40760),
            .I(N__40756));
    CascadeMux I__8759 (
            .O(N__40759),
            .I(N__40753));
    InMux I__8758 (
            .O(N__40756),
            .I(N__40748));
    InMux I__8757 (
            .O(N__40753),
            .I(N__40748));
    LocalMux I__8756 (
            .O(N__40748),
            .I(N__40744));
    InMux I__8755 (
            .O(N__40747),
            .I(N__40741));
    Span4Mux_v I__8754 (
            .O(N__40744),
            .I(N__40738));
    LocalMux I__8753 (
            .O(N__40741),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__8752 (
            .O(N__40738),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__8751 (
            .O(N__40733),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__8750 (
            .O(N__40730),
            .I(N__40726));
    CascadeMux I__8749 (
            .O(N__40729),
            .I(N__40723));
    InMux I__8748 (
            .O(N__40726),
            .I(N__40718));
    InMux I__8747 (
            .O(N__40723),
            .I(N__40718));
    LocalMux I__8746 (
            .O(N__40718),
            .I(N__40714));
    InMux I__8745 (
            .O(N__40717),
            .I(N__40711));
    Span4Mux_v I__8744 (
            .O(N__40714),
            .I(N__40708));
    LocalMux I__8743 (
            .O(N__40711),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__8742 (
            .O(N__40708),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__8741 (
            .O(N__40703),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__8740 (
            .O(N__40700),
            .I(N__40697));
    InMux I__8739 (
            .O(N__40697),
            .I(N__40694));
    LocalMux I__8738 (
            .O(N__40694),
            .I(N__40689));
    InMux I__8737 (
            .O(N__40693),
            .I(N__40686));
    InMux I__8736 (
            .O(N__40692),
            .I(N__40683));
    Span4Mux_v I__8735 (
            .O(N__40689),
            .I(N__40678));
    LocalMux I__8734 (
            .O(N__40686),
            .I(N__40678));
    LocalMux I__8733 (
            .O(N__40683),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__8732 (
            .O(N__40678),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__8731 (
            .O(N__40673),
            .I(bfn_16_23_0_));
    CascadeMux I__8730 (
            .O(N__40670),
            .I(N__40667));
    InMux I__8729 (
            .O(N__40667),
            .I(N__40664));
    LocalMux I__8728 (
            .O(N__40664),
            .I(N__40659));
    InMux I__8727 (
            .O(N__40663),
            .I(N__40656));
    InMux I__8726 (
            .O(N__40662),
            .I(N__40653));
    Span4Mux_v I__8725 (
            .O(N__40659),
            .I(N__40648));
    LocalMux I__8724 (
            .O(N__40656),
            .I(N__40648));
    LocalMux I__8723 (
            .O(N__40653),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__8722 (
            .O(N__40648),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__8721 (
            .O(N__40643),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__8720 (
            .O(N__40640),
            .I(N__40636));
    InMux I__8719 (
            .O(N__40639),
            .I(N__40633));
    LocalMux I__8718 (
            .O(N__40636),
            .I(N__40630));
    LocalMux I__8717 (
            .O(N__40633),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv4 I__8716 (
            .O(N__40630),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    CascadeMux I__8715 (
            .O(N__40625),
            .I(N__40622));
    InMux I__8714 (
            .O(N__40622),
            .I(N__40617));
    InMux I__8713 (
            .O(N__40621),
            .I(N__40614));
    InMux I__8712 (
            .O(N__40620),
            .I(N__40611));
    LocalMux I__8711 (
            .O(N__40617),
            .I(N__40606));
    LocalMux I__8710 (
            .O(N__40614),
            .I(N__40606));
    LocalMux I__8709 (
            .O(N__40611),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv4 I__8708 (
            .O(N__40606),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__8707 (
            .O(N__40601),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__8706 (
            .O(N__40598),
            .I(N__40591));
    InMux I__8705 (
            .O(N__40597),
            .I(N__40591));
    InMux I__8704 (
            .O(N__40596),
            .I(N__40588));
    LocalMux I__8703 (
            .O(N__40591),
            .I(N__40585));
    LocalMux I__8702 (
            .O(N__40588),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__8701 (
            .O(N__40585),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__8700 (
            .O(N__40580),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__8699 (
            .O(N__40577),
            .I(N__40570));
    InMux I__8698 (
            .O(N__40576),
            .I(N__40570));
    InMux I__8697 (
            .O(N__40575),
            .I(N__40567));
    LocalMux I__8696 (
            .O(N__40570),
            .I(N__40564));
    LocalMux I__8695 (
            .O(N__40567),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__8694 (
            .O(N__40564),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__8693 (
            .O(N__40559),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__8692 (
            .O(N__40556),
            .I(N__40552));
    InMux I__8691 (
            .O(N__40555),
            .I(N__40548));
    InMux I__8690 (
            .O(N__40552),
            .I(N__40545));
    InMux I__8689 (
            .O(N__40551),
            .I(N__40542));
    LocalMux I__8688 (
            .O(N__40548),
            .I(N__40537));
    LocalMux I__8687 (
            .O(N__40545),
            .I(N__40537));
    LocalMux I__8686 (
            .O(N__40542),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__8685 (
            .O(N__40537),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__8684 (
            .O(N__40532),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__8683 (
            .O(N__40529),
            .I(N__40525));
    InMux I__8682 (
            .O(N__40528),
            .I(N__40521));
    InMux I__8681 (
            .O(N__40525),
            .I(N__40518));
    InMux I__8680 (
            .O(N__40524),
            .I(N__40515));
    LocalMux I__8679 (
            .O(N__40521),
            .I(N__40510));
    LocalMux I__8678 (
            .O(N__40518),
            .I(N__40510));
    LocalMux I__8677 (
            .O(N__40515),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__8676 (
            .O(N__40510),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__8675 (
            .O(N__40505),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__8674 (
            .O(N__40502),
            .I(N__40498));
    CascadeMux I__8673 (
            .O(N__40501),
            .I(N__40495));
    InMux I__8672 (
            .O(N__40498),
            .I(N__40489));
    InMux I__8671 (
            .O(N__40495),
            .I(N__40489));
    InMux I__8670 (
            .O(N__40494),
            .I(N__40486));
    LocalMux I__8669 (
            .O(N__40489),
            .I(N__40483));
    LocalMux I__8668 (
            .O(N__40486),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__8667 (
            .O(N__40483),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__8666 (
            .O(N__40478),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__8665 (
            .O(N__40475),
            .I(N__40471));
    CascadeMux I__8664 (
            .O(N__40474),
            .I(N__40468));
    InMux I__8663 (
            .O(N__40471),
            .I(N__40462));
    InMux I__8662 (
            .O(N__40468),
            .I(N__40462));
    InMux I__8661 (
            .O(N__40467),
            .I(N__40459));
    LocalMux I__8660 (
            .O(N__40462),
            .I(N__40456));
    LocalMux I__8659 (
            .O(N__40459),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__8658 (
            .O(N__40456),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__8657 (
            .O(N__40451),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__8656 (
            .O(N__40448),
            .I(N__40445));
    InMux I__8655 (
            .O(N__40445),
            .I(N__40442));
    LocalMux I__8654 (
            .O(N__40442),
            .I(N__40437));
    InMux I__8653 (
            .O(N__40441),
            .I(N__40434));
    InMux I__8652 (
            .O(N__40440),
            .I(N__40431));
    Span4Mux_v I__8651 (
            .O(N__40437),
            .I(N__40426));
    LocalMux I__8650 (
            .O(N__40434),
            .I(N__40426));
    LocalMux I__8649 (
            .O(N__40431),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__8648 (
            .O(N__40426),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__8647 (
            .O(N__40421),
            .I(bfn_16_22_0_));
    CascadeMux I__8646 (
            .O(N__40418),
            .I(N__40415));
    InMux I__8645 (
            .O(N__40415),
            .I(N__40411));
    InMux I__8644 (
            .O(N__40414),
            .I(N__40408));
    LocalMux I__8643 (
            .O(N__40411),
            .I(N__40404));
    LocalMux I__8642 (
            .O(N__40408),
            .I(N__40401));
    InMux I__8641 (
            .O(N__40407),
            .I(N__40398));
    Span4Mux_v I__8640 (
            .O(N__40404),
            .I(N__40395));
    Span4Mux_h I__8639 (
            .O(N__40401),
            .I(N__40392));
    LocalMux I__8638 (
            .O(N__40398),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__8637 (
            .O(N__40395),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__8636 (
            .O(N__40392),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__8635 (
            .O(N__40385),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__8634 (
            .O(N__40382),
            .I(N__40379));
    InMux I__8633 (
            .O(N__40379),
            .I(N__40374));
    InMux I__8632 (
            .O(N__40378),
            .I(N__40371));
    InMux I__8631 (
            .O(N__40377),
            .I(N__40368));
    LocalMux I__8630 (
            .O(N__40374),
            .I(N__40363));
    LocalMux I__8629 (
            .O(N__40371),
            .I(N__40363));
    LocalMux I__8628 (
            .O(N__40368),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__8627 (
            .O(N__40363),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__8626 (
            .O(N__40358),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__8625 (
            .O(N__40355),
            .I(N__40348));
    InMux I__8624 (
            .O(N__40354),
            .I(N__40348));
    InMux I__8623 (
            .O(N__40353),
            .I(N__40345));
    LocalMux I__8622 (
            .O(N__40348),
            .I(N__40342));
    LocalMux I__8621 (
            .O(N__40345),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv4 I__8620 (
            .O(N__40342),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__8619 (
            .O(N__40337),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__8618 (
            .O(N__40334),
            .I(N__40330));
    CascadeMux I__8617 (
            .O(N__40333),
            .I(N__40327));
    InMux I__8616 (
            .O(N__40330),
            .I(N__40322));
    InMux I__8615 (
            .O(N__40327),
            .I(N__40322));
    LocalMux I__8614 (
            .O(N__40322),
            .I(N__40318));
    InMux I__8613 (
            .O(N__40321),
            .I(N__40315));
    Span4Mux_v I__8612 (
            .O(N__40318),
            .I(N__40312));
    LocalMux I__8611 (
            .O(N__40315),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__8610 (
            .O(N__40312),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__8609 (
            .O(N__40307),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__8608 (
            .O(N__40304),
            .I(N__40300));
    InMux I__8607 (
            .O(N__40303),
            .I(N__40296));
    InMux I__8606 (
            .O(N__40300),
            .I(N__40293));
    InMux I__8605 (
            .O(N__40299),
            .I(N__40290));
    LocalMux I__8604 (
            .O(N__40296),
            .I(N__40285));
    LocalMux I__8603 (
            .O(N__40293),
            .I(N__40285));
    LocalMux I__8602 (
            .O(N__40290),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__8601 (
            .O(N__40285),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__8600 (
            .O(N__40280),
            .I(N__40274));
    InMux I__8599 (
            .O(N__40279),
            .I(N__40271));
    InMux I__8598 (
            .O(N__40278),
            .I(N__40268));
    InMux I__8597 (
            .O(N__40277),
            .I(N__40265));
    LocalMux I__8596 (
            .O(N__40274),
            .I(N__40262));
    LocalMux I__8595 (
            .O(N__40271),
            .I(N__40259));
    LocalMux I__8594 (
            .O(N__40268),
            .I(N__40256));
    LocalMux I__8593 (
            .O(N__40265),
            .I(N__40253));
    Span4Mux_v I__8592 (
            .O(N__40262),
            .I(N__40250));
    Span4Mux_h I__8591 (
            .O(N__40259),
            .I(N__40247));
    Span4Mux_h I__8590 (
            .O(N__40256),
            .I(N__40244));
    Odrv12 I__8589 (
            .O(N__40253),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__8588 (
            .O(N__40250),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__8587 (
            .O(N__40247),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__8586 (
            .O(N__40244),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__8585 (
            .O(N__40235),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__8584 (
            .O(N__40232),
            .I(N__40225));
    InMux I__8583 (
            .O(N__40231),
            .I(N__40225));
    InMux I__8582 (
            .O(N__40230),
            .I(N__40222));
    LocalMux I__8581 (
            .O(N__40225),
            .I(N__40219));
    LocalMux I__8580 (
            .O(N__40222),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__8579 (
            .O(N__40219),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__8578 (
            .O(N__40214),
            .I(N__40208));
    InMux I__8577 (
            .O(N__40213),
            .I(N__40205));
    InMux I__8576 (
            .O(N__40212),
            .I(N__40202));
    InMux I__8575 (
            .O(N__40211),
            .I(N__40199));
    LocalMux I__8574 (
            .O(N__40208),
            .I(N__40196));
    LocalMux I__8573 (
            .O(N__40205),
            .I(N__40191));
    LocalMux I__8572 (
            .O(N__40202),
            .I(N__40191));
    LocalMux I__8571 (
            .O(N__40199),
            .I(N__40188));
    Span12Mux_h I__8570 (
            .O(N__40196),
            .I(N__40185));
    Span4Mux_v I__8569 (
            .O(N__40191),
            .I(N__40182));
    Span4Mux_h I__8568 (
            .O(N__40188),
            .I(N__40179));
    Odrv12 I__8567 (
            .O(N__40185),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__8566 (
            .O(N__40182),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__8565 (
            .O(N__40179),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__8564 (
            .O(N__40172),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__8563 (
            .O(N__40169),
            .I(N__40165));
    CascadeMux I__8562 (
            .O(N__40168),
            .I(N__40162));
    InMux I__8561 (
            .O(N__40165),
            .I(N__40156));
    InMux I__8560 (
            .O(N__40162),
            .I(N__40156));
    InMux I__8559 (
            .O(N__40161),
            .I(N__40153));
    LocalMux I__8558 (
            .O(N__40156),
            .I(N__40150));
    LocalMux I__8557 (
            .O(N__40153),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__8556 (
            .O(N__40150),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__8555 (
            .O(N__40145),
            .I(N__40141));
    InMux I__8554 (
            .O(N__40144),
            .I(N__40136));
    LocalMux I__8553 (
            .O(N__40141),
            .I(N__40133));
    InMux I__8552 (
            .O(N__40140),
            .I(N__40130));
    InMux I__8551 (
            .O(N__40139),
            .I(N__40127));
    LocalMux I__8550 (
            .O(N__40136),
            .I(N__40124));
    Span4Mux_v I__8549 (
            .O(N__40133),
            .I(N__40119));
    LocalMux I__8548 (
            .O(N__40130),
            .I(N__40119));
    LocalMux I__8547 (
            .O(N__40127),
            .I(N__40116));
    Span4Mux_h I__8546 (
            .O(N__40124),
            .I(N__40111));
    Span4Mux_h I__8545 (
            .O(N__40119),
            .I(N__40111));
    Span4Mux_h I__8544 (
            .O(N__40116),
            .I(N__40108));
    Odrv4 I__8543 (
            .O(N__40111),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__8542 (
            .O(N__40108),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__8541 (
            .O(N__40103),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__8540 (
            .O(N__40100),
            .I(N__40096));
    CascadeMux I__8539 (
            .O(N__40099),
            .I(N__40093));
    InMux I__8538 (
            .O(N__40096),
            .I(N__40087));
    InMux I__8537 (
            .O(N__40093),
            .I(N__40087));
    InMux I__8536 (
            .O(N__40092),
            .I(N__40084));
    LocalMux I__8535 (
            .O(N__40087),
            .I(N__40081));
    LocalMux I__8534 (
            .O(N__40084),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__8533 (
            .O(N__40081),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__8532 (
            .O(N__40076),
            .I(N__40071));
    InMux I__8531 (
            .O(N__40075),
            .I(N__40067));
    InMux I__8530 (
            .O(N__40074),
            .I(N__40064));
    LocalMux I__8529 (
            .O(N__40071),
            .I(N__40061));
    InMux I__8528 (
            .O(N__40070),
            .I(N__40058));
    LocalMux I__8527 (
            .O(N__40067),
            .I(N__40055));
    LocalMux I__8526 (
            .O(N__40064),
            .I(N__40052));
    Span4Mux_v I__8525 (
            .O(N__40061),
            .I(N__40049));
    LocalMux I__8524 (
            .O(N__40058),
            .I(N__40044));
    Span4Mux_v I__8523 (
            .O(N__40055),
            .I(N__40044));
    Span4Mux_h I__8522 (
            .O(N__40052),
            .I(N__40041));
    Odrv4 I__8521 (
            .O(N__40049),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    Odrv4 I__8520 (
            .O(N__40044),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    Odrv4 I__8519 (
            .O(N__40041),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__8518 (
            .O(N__40034),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__8517 (
            .O(N__40031),
            .I(N__40028));
    InMux I__8516 (
            .O(N__40028),
            .I(N__40025));
    LocalMux I__8515 (
            .O(N__40025),
            .I(N__40020));
    InMux I__8514 (
            .O(N__40024),
            .I(N__40017));
    InMux I__8513 (
            .O(N__40023),
            .I(N__40014));
    Span4Mux_v I__8512 (
            .O(N__40020),
            .I(N__40009));
    LocalMux I__8511 (
            .O(N__40017),
            .I(N__40009));
    LocalMux I__8510 (
            .O(N__40014),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__8509 (
            .O(N__40009),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__8508 (
            .O(N__40004),
            .I(N__39998));
    InMux I__8507 (
            .O(N__40003),
            .I(N__39995));
    InMux I__8506 (
            .O(N__40002),
            .I(N__39992));
    InMux I__8505 (
            .O(N__40001),
            .I(N__39989));
    LocalMux I__8504 (
            .O(N__39998),
            .I(N__39986));
    LocalMux I__8503 (
            .O(N__39995),
            .I(N__39983));
    LocalMux I__8502 (
            .O(N__39992),
            .I(N__39980));
    LocalMux I__8501 (
            .O(N__39989),
            .I(N__39977));
    Span4Mux_v I__8500 (
            .O(N__39986),
            .I(N__39972));
    Span4Mux_v I__8499 (
            .O(N__39983),
            .I(N__39972));
    Span4Mux_h I__8498 (
            .O(N__39980),
            .I(N__39967));
    Span4Mux_h I__8497 (
            .O(N__39977),
            .I(N__39967));
    Odrv4 I__8496 (
            .O(N__39972),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    Odrv4 I__8495 (
            .O(N__39967),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__8494 (
            .O(N__39962),
            .I(bfn_16_21_0_));
    CascadeMux I__8493 (
            .O(N__39959),
            .I(N__39956));
    InMux I__8492 (
            .O(N__39956),
            .I(N__39953));
    LocalMux I__8491 (
            .O(N__39953),
            .I(N__39948));
    InMux I__8490 (
            .O(N__39952),
            .I(N__39945));
    InMux I__8489 (
            .O(N__39951),
            .I(N__39942));
    Span4Mux_v I__8488 (
            .O(N__39948),
            .I(N__39937));
    LocalMux I__8487 (
            .O(N__39945),
            .I(N__39937));
    LocalMux I__8486 (
            .O(N__39942),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__8485 (
            .O(N__39937),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__8484 (
            .O(N__39932),
            .I(N__39929));
    LocalMux I__8483 (
            .O(N__39929),
            .I(N__39924));
    InMux I__8482 (
            .O(N__39928),
            .I(N__39921));
    InMux I__8481 (
            .O(N__39927),
            .I(N__39917));
    Span4Mux_h I__8480 (
            .O(N__39924),
            .I(N__39912));
    LocalMux I__8479 (
            .O(N__39921),
            .I(N__39912));
    CascadeMux I__8478 (
            .O(N__39920),
            .I(N__39909));
    LocalMux I__8477 (
            .O(N__39917),
            .I(N__39906));
    Span4Mux_h I__8476 (
            .O(N__39912),
            .I(N__39903));
    InMux I__8475 (
            .O(N__39909),
            .I(N__39900));
    Span4Mux_h I__8474 (
            .O(N__39906),
            .I(N__39895));
    Span4Mux_v I__8473 (
            .O(N__39903),
            .I(N__39895));
    LocalMux I__8472 (
            .O(N__39900),
            .I(N__39892));
    Span4Mux_v I__8471 (
            .O(N__39895),
            .I(N__39889));
    Span4Mux_h I__8470 (
            .O(N__39892),
            .I(N__39886));
    Odrv4 I__8469 (
            .O(N__39889),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__8468 (
            .O(N__39886),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__8467 (
            .O(N__39881),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__8466 (
            .O(N__39878),
            .I(N__39875));
    LocalMux I__8465 (
            .O(N__39875),
            .I(N__39870));
    InMux I__8464 (
            .O(N__39874),
            .I(N__39865));
    InMux I__8463 (
            .O(N__39873),
            .I(N__39865));
    Odrv4 I__8462 (
            .O(N__39870),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__8461 (
            .O(N__39865),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    InMux I__8460 (
            .O(N__39860),
            .I(N__39857));
    LocalMux I__8459 (
            .O(N__39857),
            .I(N__39853));
    InMux I__8458 (
            .O(N__39856),
            .I(N__39850));
    Span4Mux_h I__8457 (
            .O(N__39853),
            .I(N__39847));
    LocalMux I__8456 (
            .O(N__39850),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    Odrv4 I__8455 (
            .O(N__39847),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    CascadeMux I__8454 (
            .O(N__39842),
            .I(elapsed_time_ns_1_RNI14DN9_0_23_cascade_));
    InMux I__8453 (
            .O(N__39839),
            .I(N__39833));
    InMux I__8452 (
            .O(N__39838),
            .I(N__39833));
    LocalMux I__8451 (
            .O(N__39833),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    InMux I__8450 (
            .O(N__39830),
            .I(N__39827));
    LocalMux I__8449 (
            .O(N__39827),
            .I(N__39824));
    Span4Mux_v I__8448 (
            .O(N__39824),
            .I(N__39820));
    InMux I__8447 (
            .O(N__39823),
            .I(N__39817));
    Odrv4 I__8446 (
            .O(N__39820),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    LocalMux I__8445 (
            .O(N__39817),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    CascadeMux I__8444 (
            .O(N__39812),
            .I(elapsed_time_ns_1_RNI03DN9_0_22_cascade_));
    InMux I__8443 (
            .O(N__39809),
            .I(N__39803));
    InMux I__8442 (
            .O(N__39808),
            .I(N__39803));
    LocalMux I__8441 (
            .O(N__39803),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ));
    CascadeMux I__8440 (
            .O(N__39800),
            .I(N__39796));
    InMux I__8439 (
            .O(N__39799),
            .I(N__39793));
    InMux I__8438 (
            .O(N__39796),
            .I(N__39790));
    LocalMux I__8437 (
            .O(N__39793),
            .I(N__39784));
    LocalMux I__8436 (
            .O(N__39790),
            .I(N__39784));
    InMux I__8435 (
            .O(N__39789),
            .I(N__39781));
    Span4Mux_v I__8434 (
            .O(N__39784),
            .I(N__39778));
    LocalMux I__8433 (
            .O(N__39781),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv4 I__8432 (
            .O(N__39778),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__8431 (
            .O(N__39773),
            .I(N__39768));
    InMux I__8430 (
            .O(N__39772),
            .I(N__39765));
    CascadeMux I__8429 (
            .O(N__39771),
            .I(N__39761));
    LocalMux I__8428 (
            .O(N__39768),
            .I(N__39758));
    LocalMux I__8427 (
            .O(N__39765),
            .I(N__39755));
    InMux I__8426 (
            .O(N__39764),
            .I(N__39750));
    InMux I__8425 (
            .O(N__39761),
            .I(N__39750));
    Span4Mux_v I__8424 (
            .O(N__39758),
            .I(N__39743));
    Span4Mux_v I__8423 (
            .O(N__39755),
            .I(N__39743));
    LocalMux I__8422 (
            .O(N__39750),
            .I(N__39743));
    Odrv4 I__8421 (
            .O(N__39743),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__8420 (
            .O(N__39740),
            .I(N__39736));
    InMux I__8419 (
            .O(N__39739),
            .I(N__39733));
    LocalMux I__8418 (
            .O(N__39736),
            .I(N__39727));
    LocalMux I__8417 (
            .O(N__39733),
            .I(N__39727));
    InMux I__8416 (
            .O(N__39732),
            .I(N__39724));
    Span4Mux_v I__8415 (
            .O(N__39727),
            .I(N__39721));
    LocalMux I__8414 (
            .O(N__39724),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__8413 (
            .O(N__39721),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__8412 (
            .O(N__39716),
            .I(N__39712));
    InMux I__8411 (
            .O(N__39715),
            .I(N__39707));
    LocalMux I__8410 (
            .O(N__39712),
            .I(N__39704));
    InMux I__8409 (
            .O(N__39711),
            .I(N__39699));
    InMux I__8408 (
            .O(N__39710),
            .I(N__39699));
    LocalMux I__8407 (
            .O(N__39707),
            .I(N__39696));
    Span4Mux_v I__8406 (
            .O(N__39704),
            .I(N__39691));
    LocalMux I__8405 (
            .O(N__39699),
            .I(N__39691));
    Odrv12 I__8404 (
            .O(N__39696),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__8403 (
            .O(N__39691),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__8402 (
            .O(N__39686),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__8401 (
            .O(N__39683),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ));
    InMux I__8400 (
            .O(N__39680),
            .I(N__39674));
    InMux I__8399 (
            .O(N__39679),
            .I(N__39674));
    LocalMux I__8398 (
            .O(N__39674),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    CascadeMux I__8397 (
            .O(N__39671),
            .I(N__39666));
    InMux I__8396 (
            .O(N__39670),
            .I(N__39660));
    InMux I__8395 (
            .O(N__39669),
            .I(N__39660));
    InMux I__8394 (
            .O(N__39666),
            .I(N__39655));
    InMux I__8393 (
            .O(N__39665),
            .I(N__39655));
    LocalMux I__8392 (
            .O(N__39660),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__8391 (
            .O(N__39655),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    InMux I__8390 (
            .O(N__39650),
            .I(N__39641));
    InMux I__8389 (
            .O(N__39649),
            .I(N__39641));
    InMux I__8388 (
            .O(N__39648),
            .I(N__39641));
    LocalMux I__8387 (
            .O(N__39641),
            .I(N__39638));
    Odrv4 I__8386 (
            .O(N__39638),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    InMux I__8385 (
            .O(N__39635),
            .I(N__39626));
    InMux I__8384 (
            .O(N__39634),
            .I(N__39626));
    InMux I__8383 (
            .O(N__39633),
            .I(N__39626));
    LocalMux I__8382 (
            .O(N__39626),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    CascadeMux I__8381 (
            .O(N__39623),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ));
    InMux I__8380 (
            .O(N__39620),
            .I(N__39617));
    LocalMux I__8379 (
            .O(N__39617),
            .I(N__39614));
    Odrv4 I__8378 (
            .O(N__39614),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__8377 (
            .O(N__39611),
            .I(N__39607));
    InMux I__8376 (
            .O(N__39610),
            .I(N__39604));
    LocalMux I__8375 (
            .O(N__39607),
            .I(N__39601));
    LocalMux I__8374 (
            .O(N__39604),
            .I(N__39598));
    Span4Mux_h I__8373 (
            .O(N__39601),
            .I(N__39595));
    Span4Mux_h I__8372 (
            .O(N__39598),
            .I(N__39588));
    Span4Mux_v I__8371 (
            .O(N__39595),
            .I(N__39588));
    InMux I__8370 (
            .O(N__39594),
            .I(N__39583));
    InMux I__8369 (
            .O(N__39593),
            .I(N__39583));
    Span4Mux_v I__8368 (
            .O(N__39588),
            .I(N__39580));
    LocalMux I__8367 (
            .O(N__39583),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__8366 (
            .O(N__39580),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    CEMux I__8365 (
            .O(N__39575),
            .I(N__39571));
    CEMux I__8364 (
            .O(N__39574),
            .I(N__39566));
    LocalMux I__8363 (
            .O(N__39571),
            .I(N__39563));
    CEMux I__8362 (
            .O(N__39570),
            .I(N__39560));
    CEMux I__8361 (
            .O(N__39569),
            .I(N__39557));
    LocalMux I__8360 (
            .O(N__39566),
            .I(N__39554));
    Span4Mux_v I__8359 (
            .O(N__39563),
            .I(N__39547));
    LocalMux I__8358 (
            .O(N__39560),
            .I(N__39547));
    LocalMux I__8357 (
            .O(N__39557),
            .I(N__39547));
    Span4Mux_v I__8356 (
            .O(N__39554),
            .I(N__39542));
    Span4Mux_v I__8355 (
            .O(N__39547),
            .I(N__39542));
    Odrv4 I__8354 (
            .O(N__39542),
            .I(\delay_measurement_inst.delay_hc_timer.N_202_i ));
    InMux I__8353 (
            .O(N__39539),
            .I(N__39525));
    InMux I__8352 (
            .O(N__39538),
            .I(N__39525));
    InMux I__8351 (
            .O(N__39537),
            .I(N__39525));
    InMux I__8350 (
            .O(N__39536),
            .I(N__39525));
    InMux I__8349 (
            .O(N__39535),
            .I(N__39496));
    InMux I__8348 (
            .O(N__39534),
            .I(N__39496));
    LocalMux I__8347 (
            .O(N__39525),
            .I(N__39493));
    InMux I__8346 (
            .O(N__39524),
            .I(N__39484));
    InMux I__8345 (
            .O(N__39523),
            .I(N__39484));
    InMux I__8344 (
            .O(N__39522),
            .I(N__39484));
    InMux I__8343 (
            .O(N__39521),
            .I(N__39484));
    InMux I__8342 (
            .O(N__39520),
            .I(N__39475));
    InMux I__8341 (
            .O(N__39519),
            .I(N__39475));
    InMux I__8340 (
            .O(N__39518),
            .I(N__39475));
    InMux I__8339 (
            .O(N__39517),
            .I(N__39475));
    InMux I__8338 (
            .O(N__39516),
            .I(N__39466));
    InMux I__8337 (
            .O(N__39515),
            .I(N__39466));
    InMux I__8336 (
            .O(N__39514),
            .I(N__39466));
    InMux I__8335 (
            .O(N__39513),
            .I(N__39466));
    InMux I__8334 (
            .O(N__39512),
            .I(N__39457));
    InMux I__8333 (
            .O(N__39511),
            .I(N__39457));
    InMux I__8332 (
            .O(N__39510),
            .I(N__39457));
    InMux I__8331 (
            .O(N__39509),
            .I(N__39457));
    InMux I__8330 (
            .O(N__39508),
            .I(N__39448));
    InMux I__8329 (
            .O(N__39507),
            .I(N__39448));
    InMux I__8328 (
            .O(N__39506),
            .I(N__39448));
    InMux I__8327 (
            .O(N__39505),
            .I(N__39448));
    InMux I__8326 (
            .O(N__39504),
            .I(N__39439));
    InMux I__8325 (
            .O(N__39503),
            .I(N__39439));
    InMux I__8324 (
            .O(N__39502),
            .I(N__39439));
    InMux I__8323 (
            .O(N__39501),
            .I(N__39439));
    LocalMux I__8322 (
            .O(N__39496),
            .I(N__39436));
    Span4Mux_h I__8321 (
            .O(N__39493),
            .I(N__39431));
    LocalMux I__8320 (
            .O(N__39484),
            .I(N__39431));
    LocalMux I__8319 (
            .O(N__39475),
            .I(N__39418));
    LocalMux I__8318 (
            .O(N__39466),
            .I(N__39418));
    LocalMux I__8317 (
            .O(N__39457),
            .I(N__39418));
    LocalMux I__8316 (
            .O(N__39448),
            .I(N__39418));
    LocalMux I__8315 (
            .O(N__39439),
            .I(N__39418));
    Span4Mux_h I__8314 (
            .O(N__39436),
            .I(N__39418));
    Span4Mux_v I__8313 (
            .O(N__39431),
            .I(N__39415));
    Span4Mux_v I__8312 (
            .O(N__39418),
            .I(N__39412));
    Odrv4 I__8311 (
            .O(N__39415),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__8310 (
            .O(N__39412),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__8309 (
            .O(N__39407),
            .I(N__39402));
    InMux I__8308 (
            .O(N__39406),
            .I(N__39397));
    InMux I__8307 (
            .O(N__39405),
            .I(N__39397));
    LocalMux I__8306 (
            .O(N__39402),
            .I(N__39391));
    LocalMux I__8305 (
            .O(N__39397),
            .I(N__39391));
    InMux I__8304 (
            .O(N__39396),
            .I(N__39388));
    Span12Mux_v I__8303 (
            .O(N__39391),
            .I(N__39385));
    LocalMux I__8302 (
            .O(N__39388),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__8301 (
            .O(N__39385),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__8300 (
            .O(N__39380),
            .I(N__39376));
    InMux I__8299 (
            .O(N__39379),
            .I(N__39372));
    LocalMux I__8298 (
            .O(N__39376),
            .I(N__39369));
    InMux I__8297 (
            .O(N__39375),
            .I(N__39366));
    LocalMux I__8296 (
            .O(N__39372),
            .I(N__39363));
    Span4Mux_h I__8295 (
            .O(N__39369),
            .I(N__39360));
    LocalMux I__8294 (
            .O(N__39366),
            .I(N__39357));
    Span4Mux_h I__8293 (
            .O(N__39363),
            .I(N__39352));
    Span4Mux_v I__8292 (
            .O(N__39360),
            .I(N__39352));
    Span4Mux_h I__8291 (
            .O(N__39357),
            .I(N__39349));
    Span4Mux_v I__8290 (
            .O(N__39352),
            .I(N__39346));
    Sp12to4 I__8289 (
            .O(N__39349),
            .I(N__39343));
    Odrv4 I__8288 (
            .O(N__39346),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv12 I__8287 (
            .O(N__39343),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__8286 (
            .O(N__39338),
            .I(N__39335));
    LocalMux I__8285 (
            .O(N__39335),
            .I(N__39331));
    InMux I__8284 (
            .O(N__39334),
            .I(N__39327));
    Span4Mux_v I__8283 (
            .O(N__39331),
            .I(N__39324));
    InMux I__8282 (
            .O(N__39330),
            .I(N__39321));
    LocalMux I__8281 (
            .O(N__39327),
            .I(N__39318));
    Span4Mux_v I__8280 (
            .O(N__39324),
            .I(N__39315));
    LocalMux I__8279 (
            .O(N__39321),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv4 I__8278 (
            .O(N__39318),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv4 I__8277 (
            .O(N__39315),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    InMux I__8276 (
            .O(N__39308),
            .I(N__39304));
    InMux I__8275 (
            .O(N__39307),
            .I(N__39300));
    LocalMux I__8274 (
            .O(N__39304),
            .I(N__39297));
    InMux I__8273 (
            .O(N__39303),
            .I(N__39294));
    LocalMux I__8272 (
            .O(N__39300),
            .I(N__39291));
    Span12Mux_v I__8271 (
            .O(N__39297),
            .I(N__39288));
    LocalMux I__8270 (
            .O(N__39294),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    Odrv4 I__8269 (
            .O(N__39291),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    Odrv12 I__8268 (
            .O(N__39288),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    InMux I__8267 (
            .O(N__39281),
            .I(N__39276));
    InMux I__8266 (
            .O(N__39280),
            .I(N__39273));
    InMux I__8265 (
            .O(N__39279),
            .I(N__39270));
    LocalMux I__8264 (
            .O(N__39276),
            .I(N__39267));
    LocalMux I__8263 (
            .O(N__39273),
            .I(N__39264));
    LocalMux I__8262 (
            .O(N__39270),
            .I(N__39259));
    Span4Mux_v I__8261 (
            .O(N__39267),
            .I(N__39259));
    Odrv12 I__8260 (
            .O(N__39264),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    Odrv4 I__8259 (
            .O(N__39259),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    InMux I__8258 (
            .O(N__39254),
            .I(N__39248));
    InMux I__8257 (
            .O(N__39253),
            .I(N__39243));
    InMux I__8256 (
            .O(N__39252),
            .I(N__39243));
    InMux I__8255 (
            .O(N__39251),
            .I(N__39240));
    LocalMux I__8254 (
            .O(N__39248),
            .I(N__39235));
    LocalMux I__8253 (
            .O(N__39243),
            .I(N__39235));
    LocalMux I__8252 (
            .O(N__39240),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv12 I__8251 (
            .O(N__39235),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__8250 (
            .O(N__39230),
            .I(N__39220));
    InMux I__8249 (
            .O(N__39229),
            .I(N__39220));
    InMux I__8248 (
            .O(N__39228),
            .I(N__39220));
    InMux I__8247 (
            .O(N__39227),
            .I(N__39216));
    LocalMux I__8246 (
            .O(N__39220),
            .I(N__39211));
    InMux I__8245 (
            .O(N__39219),
            .I(N__39208));
    LocalMux I__8244 (
            .O(N__39216),
            .I(N__39205));
    InMux I__8243 (
            .O(N__39215),
            .I(N__39202));
    InMux I__8242 (
            .O(N__39214),
            .I(N__39199));
    Span4Mux_v I__8241 (
            .O(N__39211),
            .I(N__39196));
    LocalMux I__8240 (
            .O(N__39208),
            .I(N__39188));
    Span4Mux_h I__8239 (
            .O(N__39205),
            .I(N__39188));
    LocalMux I__8238 (
            .O(N__39202),
            .I(N__39188));
    LocalMux I__8237 (
            .O(N__39199),
            .I(N__39183));
    Span4Mux_v I__8236 (
            .O(N__39196),
            .I(N__39183));
    InMux I__8235 (
            .O(N__39195),
            .I(N__39180));
    Odrv4 I__8234 (
            .O(N__39188),
            .I(state_3));
    Odrv4 I__8233 (
            .O(N__39183),
            .I(state_3));
    LocalMux I__8232 (
            .O(N__39180),
            .I(state_3));
    InMux I__8231 (
            .O(N__39173),
            .I(N__39169));
    InMux I__8230 (
            .O(N__39172),
            .I(N__39163));
    LocalMux I__8229 (
            .O(N__39169),
            .I(N__39160));
    InMux I__8228 (
            .O(N__39168),
            .I(N__39157));
    InMux I__8227 (
            .O(N__39167),
            .I(N__39152));
    InMux I__8226 (
            .O(N__39166),
            .I(N__39152));
    LocalMux I__8225 (
            .O(N__39163),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__8224 (
            .O(N__39160),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__8223 (
            .O(N__39157),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__8222 (
            .O(N__39152),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    IoInMux I__8221 (
            .O(N__39143),
            .I(N__39140));
    LocalMux I__8220 (
            .O(N__39140),
            .I(N__39137));
    Span4Mux_s2_v I__8219 (
            .O(N__39137),
            .I(N__39134));
    Span4Mux_v I__8218 (
            .O(N__39134),
            .I(N__39131));
    Span4Mux_v I__8217 (
            .O(N__39131),
            .I(N__39128));
    Span4Mux_v I__8216 (
            .O(N__39128),
            .I(N__39124));
    InMux I__8215 (
            .O(N__39127),
            .I(N__39121));
    Odrv4 I__8214 (
            .O(N__39124),
            .I(T01_c));
    LocalMux I__8213 (
            .O(N__39121),
            .I(T01_c));
    InMux I__8212 (
            .O(N__39116),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__8211 (
            .O(N__39113),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__8210 (
            .O(N__39110),
            .I(N__39107));
    LocalMux I__8209 (
            .O(N__39107),
            .I(N__39103));
    InMux I__8208 (
            .O(N__39106),
            .I(N__39099));
    Span4Mux_v I__8207 (
            .O(N__39103),
            .I(N__39096));
    InMux I__8206 (
            .O(N__39102),
            .I(N__39093));
    LocalMux I__8205 (
            .O(N__39099),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__8204 (
            .O(N__39096),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__8203 (
            .O(N__39093),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__8202 (
            .O(N__39086),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__8201 (
            .O(N__39083),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__8200 (
            .O(N__39080),
            .I(N__39076));
    CascadeMux I__8199 (
            .O(N__39079),
            .I(N__39072));
    InMux I__8198 (
            .O(N__39076),
            .I(N__39067));
    InMux I__8197 (
            .O(N__39075),
            .I(N__39067));
    InMux I__8196 (
            .O(N__39072),
            .I(N__39064));
    LocalMux I__8195 (
            .O(N__39067),
            .I(N__39061));
    LocalMux I__8194 (
            .O(N__39064),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv4 I__8193 (
            .O(N__39061),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    InMux I__8192 (
            .O(N__39056),
            .I(N__39053));
    LocalMux I__8191 (
            .O(N__39053),
            .I(N__39050));
    Odrv4 I__8190 (
            .O(N__39050),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    CascadeMux I__8189 (
            .O(N__39047),
            .I(N__39044));
    InMux I__8188 (
            .O(N__39044),
            .I(N__39041));
    LocalMux I__8187 (
            .O(N__39041),
            .I(N__39038));
    Span4Mux_h I__8186 (
            .O(N__39038),
            .I(N__39035));
    Span4Mux_v I__8185 (
            .O(N__39035),
            .I(N__39032));
    Odrv4 I__8184 (
            .O(N__39032),
            .I(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ));
    InMux I__8183 (
            .O(N__39029),
            .I(N__39026));
    LocalMux I__8182 (
            .O(N__39026),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__8181 (
            .O(N__39023),
            .I(N__39020));
    LocalMux I__8180 (
            .O(N__39020),
            .I(N__39017));
    Odrv4 I__8179 (
            .O(N__39017),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    CascadeMux I__8178 (
            .O(N__39014),
            .I(N__39011));
    InMux I__8177 (
            .O(N__39011),
            .I(N__39008));
    LocalMux I__8176 (
            .O(N__39008),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__8175 (
            .O(N__39005),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__8174 (
            .O(N__39002),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__8173 (
            .O(N__38999),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__8172 (
            .O(N__38996),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__8171 (
            .O(N__38993),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__8170 (
            .O(N__38990),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    CascadeMux I__8169 (
            .O(N__38987),
            .I(N__38984));
    InMux I__8168 (
            .O(N__38984),
            .I(N__38981));
    LocalMux I__8167 (
            .O(N__38981),
            .I(N__38977));
    InMux I__8166 (
            .O(N__38980),
            .I(N__38974));
    Span4Mux_v I__8165 (
            .O(N__38977),
            .I(N__38968));
    LocalMux I__8164 (
            .O(N__38974),
            .I(N__38968));
    InMux I__8163 (
            .O(N__38973),
            .I(N__38965));
    Span4Mux_h I__8162 (
            .O(N__38968),
            .I(N__38962));
    LocalMux I__8161 (
            .O(N__38965),
            .I(N__38959));
    Odrv4 I__8160 (
            .O(N__38962),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv12 I__8159 (
            .O(N__38959),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__8158 (
            .O(N__38954),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__8157 (
            .O(N__38951),
            .I(bfn_16_11_0_));
    InMux I__8156 (
            .O(N__38948),
            .I(N__38945));
    LocalMux I__8155 (
            .O(N__38945),
            .I(N__38942));
    Span4Mux_h I__8154 (
            .O(N__38942),
            .I(N__38937));
    InMux I__8153 (
            .O(N__38941),
            .I(N__38932));
    InMux I__8152 (
            .O(N__38940),
            .I(N__38932));
    Odrv4 I__8151 (
            .O(N__38937),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__8150 (
            .O(N__38932),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__8149 (
            .O(N__38927),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__8148 (
            .O(N__38924),
            .I(N__38921));
    LocalMux I__8147 (
            .O(N__38921),
            .I(N__38918));
    Span4Mux_v I__8146 (
            .O(N__38918),
            .I(N__38915));
    Odrv4 I__8145 (
            .O(N__38915),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    CascadeMux I__8144 (
            .O(N__38912),
            .I(N__38908));
    InMux I__8143 (
            .O(N__38911),
            .I(N__38905));
    InMux I__8142 (
            .O(N__38908),
            .I(N__38901));
    LocalMux I__8141 (
            .O(N__38905),
            .I(N__38898));
    InMux I__8140 (
            .O(N__38904),
            .I(N__38895));
    LocalMux I__8139 (
            .O(N__38901),
            .I(N__38892));
    Span4Mux_h I__8138 (
            .O(N__38898),
            .I(N__38889));
    LocalMux I__8137 (
            .O(N__38895),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv4 I__8136 (
            .O(N__38892),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv4 I__8135 (
            .O(N__38889),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__8134 (
            .O(N__38882),
            .I(bfn_16_9_0_));
    InMux I__8133 (
            .O(N__38879),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__8132 (
            .O(N__38876),
            .I(N__38873));
    LocalMux I__8131 (
            .O(N__38873),
            .I(N__38868));
    InMux I__8130 (
            .O(N__38872),
            .I(N__38865));
    InMux I__8129 (
            .O(N__38871),
            .I(N__38862));
    Odrv4 I__8128 (
            .O(N__38868),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__8127 (
            .O(N__38865),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__8126 (
            .O(N__38862),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__8125 (
            .O(N__38855),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__8124 (
            .O(N__38852),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__8123 (
            .O(N__38849),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__8122 (
            .O(N__38846),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__8121 (
            .O(N__38843),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__8120 (
            .O(N__38840),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__8119 (
            .O(N__38837),
            .I(bfn_16_10_0_));
    InMux I__8118 (
            .O(N__38834),
            .I(N__38831));
    LocalMux I__8117 (
            .O(N__38831),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    InMux I__8116 (
            .O(N__38828),
            .I(N__38823));
    CascadeMux I__8115 (
            .O(N__38827),
            .I(N__38820));
    InMux I__8114 (
            .O(N__38826),
            .I(N__38817));
    LocalMux I__8113 (
            .O(N__38823),
            .I(N__38814));
    InMux I__8112 (
            .O(N__38820),
            .I(N__38811));
    LocalMux I__8111 (
            .O(N__38817),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__8110 (
            .O(N__38814),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__8109 (
            .O(N__38811),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__8108 (
            .O(N__38804),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__8107 (
            .O(N__38801),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__8106 (
            .O(N__38798),
            .I(N__38795));
    LocalMux I__8105 (
            .O(N__38795),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__8104 (
            .O(N__38792),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__8103 (
            .O(N__38789),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__8102 (
            .O(N__38786),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__8101 (
            .O(N__38783),
            .I(N__38780));
    LocalMux I__8100 (
            .O(N__38780),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__8099 (
            .O(N__38777),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__8098 (
            .O(N__38774),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__8097 (
            .O(N__38771),
            .I(N__38768));
    LocalMux I__8096 (
            .O(N__38768),
            .I(N__38765));
    Odrv4 I__8095 (
            .O(N__38765),
            .I(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ));
    CascadeMux I__8094 (
            .O(N__38762),
            .I(N__38759));
    InMux I__8093 (
            .O(N__38759),
            .I(N__38756));
    LocalMux I__8092 (
            .O(N__38756),
            .I(N__38753));
    Odrv4 I__8091 (
            .O(N__38753),
            .I(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ));
    CascadeMux I__8090 (
            .O(N__38750),
            .I(N__38747));
    InMux I__8089 (
            .O(N__38747),
            .I(N__38744));
    LocalMux I__8088 (
            .O(N__38744),
            .I(N__38741));
    Odrv12 I__8087 (
            .O(N__38741),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    CascadeMux I__8086 (
            .O(N__38738),
            .I(N__38735));
    InMux I__8085 (
            .O(N__38735),
            .I(N__38732));
    LocalMux I__8084 (
            .O(N__38732),
            .I(N__38729));
    Odrv12 I__8083 (
            .O(N__38729),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    CascadeMux I__8082 (
            .O(N__38726),
            .I(N__38723));
    InMux I__8081 (
            .O(N__38723),
            .I(N__38720));
    LocalMux I__8080 (
            .O(N__38720),
            .I(N__38717));
    Odrv4 I__8079 (
            .O(N__38717),
            .I(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ));
    CascadeMux I__8078 (
            .O(N__38714),
            .I(N__38711));
    InMux I__8077 (
            .O(N__38711),
            .I(N__38708));
    LocalMux I__8076 (
            .O(N__38708),
            .I(N__38705));
    Span4Mux_h I__8075 (
            .O(N__38705),
            .I(N__38702));
    Odrv4 I__8074 (
            .O(N__38702),
            .I(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ));
    CascadeMux I__8073 (
            .O(N__38699),
            .I(N__38696));
    InMux I__8072 (
            .O(N__38696),
            .I(N__38693));
    LocalMux I__8071 (
            .O(N__38693),
            .I(N__38690));
    Sp12to4 I__8070 (
            .O(N__38690),
            .I(N__38687));
    Odrv12 I__8069 (
            .O(N__38687),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    CascadeMux I__8068 (
            .O(N__38684),
            .I(N__38681));
    InMux I__8067 (
            .O(N__38681),
            .I(N__38678));
    LocalMux I__8066 (
            .O(N__38678),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    CascadeMux I__8065 (
            .O(N__38675),
            .I(N__38671));
    InMux I__8064 (
            .O(N__38674),
            .I(N__38666));
    InMux I__8063 (
            .O(N__38671),
            .I(N__38666));
    LocalMux I__8062 (
            .O(N__38666),
            .I(N__38662));
    InMux I__8061 (
            .O(N__38665),
            .I(N__38659));
    Span4Mux_v I__8060 (
            .O(N__38662),
            .I(N__38656));
    LocalMux I__8059 (
            .O(N__38659),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__8058 (
            .O(N__38656),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__8057 (
            .O(N__38651),
            .I(N__38647));
    InMux I__8056 (
            .O(N__38650),
            .I(N__38642));
    InMux I__8055 (
            .O(N__38647),
            .I(N__38642));
    LocalMux I__8054 (
            .O(N__38642),
            .I(N__38638));
    InMux I__8053 (
            .O(N__38641),
            .I(N__38635));
    Span4Mux_v I__8052 (
            .O(N__38638),
            .I(N__38632));
    LocalMux I__8051 (
            .O(N__38635),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__8050 (
            .O(N__38632),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__8049 (
            .O(N__38627),
            .I(N__38621));
    InMux I__8048 (
            .O(N__38626),
            .I(N__38621));
    LocalMux I__8047 (
            .O(N__38621),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__8046 (
            .O(N__38618),
            .I(N__38615));
    LocalMux I__8045 (
            .O(N__38615),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    InMux I__8044 (
            .O(N__38612),
            .I(N__38609));
    LocalMux I__8043 (
            .O(N__38609),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    InMux I__8042 (
            .O(N__38606),
            .I(N__38603));
    LocalMux I__8041 (
            .O(N__38603),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    CascadeMux I__8040 (
            .O(N__38600),
            .I(N__38596));
    CascadeMux I__8039 (
            .O(N__38599),
            .I(N__38593));
    InMux I__8038 (
            .O(N__38596),
            .I(N__38589));
    InMux I__8037 (
            .O(N__38593),
            .I(N__38586));
    InMux I__8036 (
            .O(N__38592),
            .I(N__38583));
    LocalMux I__8035 (
            .O(N__38589),
            .I(N__38579));
    LocalMux I__8034 (
            .O(N__38586),
            .I(N__38574));
    LocalMux I__8033 (
            .O(N__38583),
            .I(N__38574));
    InMux I__8032 (
            .O(N__38582),
            .I(N__38571));
    Span4Mux_v I__8031 (
            .O(N__38579),
            .I(N__38568));
    Span4Mux_v I__8030 (
            .O(N__38574),
            .I(N__38565));
    LocalMux I__8029 (
            .O(N__38571),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__8028 (
            .O(N__38568),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__8027 (
            .O(N__38565),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__8026 (
            .O(N__38558),
            .I(N__38554));
    InMux I__8025 (
            .O(N__38557),
            .I(N__38550));
    InMux I__8024 (
            .O(N__38554),
            .I(N__38547));
    InMux I__8023 (
            .O(N__38553),
            .I(N__38544));
    LocalMux I__8022 (
            .O(N__38550),
            .I(N__38538));
    LocalMux I__8021 (
            .O(N__38547),
            .I(N__38538));
    LocalMux I__8020 (
            .O(N__38544),
            .I(N__38535));
    InMux I__8019 (
            .O(N__38543),
            .I(N__38532));
    Span4Mux_v I__8018 (
            .O(N__38538),
            .I(N__38529));
    Span4Mux_v I__8017 (
            .O(N__38535),
            .I(N__38526));
    LocalMux I__8016 (
            .O(N__38532),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__8015 (
            .O(N__38529),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__8014 (
            .O(N__38526),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    CascadeMux I__8013 (
            .O(N__38519),
            .I(N__38516));
    InMux I__8012 (
            .O(N__38516),
            .I(N__38512));
    InMux I__8011 (
            .O(N__38515),
            .I(N__38509));
    LocalMux I__8010 (
            .O(N__38512),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    LocalMux I__8009 (
            .O(N__38509),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    InMux I__8008 (
            .O(N__38504),
            .I(N__38501));
    LocalMux I__8007 (
            .O(N__38501),
            .I(N__38498));
    Span4Mux_v I__8006 (
            .O(N__38498),
            .I(N__38495));
    Odrv4 I__8005 (
            .O(N__38495),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    InMux I__8004 (
            .O(N__38492),
            .I(N__38489));
    LocalMux I__8003 (
            .O(N__38489),
            .I(N__38486));
    Odrv4 I__8002 (
            .O(N__38486),
            .I(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ));
    InMux I__8001 (
            .O(N__38483),
            .I(N__38480));
    LocalMux I__8000 (
            .O(N__38480),
            .I(N__38477));
    Odrv12 I__7999 (
            .O(N__38477),
            .I(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ));
    InMux I__7998 (
            .O(N__38474),
            .I(N__38469));
    InMux I__7997 (
            .O(N__38473),
            .I(N__38466));
    InMux I__7996 (
            .O(N__38472),
            .I(N__38463));
    LocalMux I__7995 (
            .O(N__38469),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__7994 (
            .O(N__38466),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__7993 (
            .O(N__38463),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    CascadeMux I__7992 (
            .O(N__38456),
            .I(N__38452));
    CascadeMux I__7991 (
            .O(N__38455),
            .I(N__38448));
    InMux I__7990 (
            .O(N__38452),
            .I(N__38445));
    InMux I__7989 (
            .O(N__38451),
            .I(N__38442));
    InMux I__7988 (
            .O(N__38448),
            .I(N__38439));
    LocalMux I__7987 (
            .O(N__38445),
            .I(N__38436));
    LocalMux I__7986 (
            .O(N__38442),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__7985 (
            .O(N__38439),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv4 I__7984 (
            .O(N__38436),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    CascadeMux I__7983 (
            .O(N__38429),
            .I(N__38426));
    InMux I__7982 (
            .O(N__38426),
            .I(N__38423));
    LocalMux I__7981 (
            .O(N__38423),
            .I(N__38420));
    Span4Mux_v I__7980 (
            .O(N__38420),
            .I(N__38417));
    Odrv4 I__7979 (
            .O(N__38417),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt26 ));
    InMux I__7978 (
            .O(N__38414),
            .I(N__38411));
    LocalMux I__7977 (
            .O(N__38411),
            .I(N__38408));
    Odrv4 I__7976 (
            .O(N__38408),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ));
    InMux I__7975 (
            .O(N__38405),
            .I(N__38400));
    InMux I__7974 (
            .O(N__38404),
            .I(N__38395));
    InMux I__7973 (
            .O(N__38403),
            .I(N__38395));
    LocalMux I__7972 (
            .O(N__38400),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__7971 (
            .O(N__38395),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    CascadeMux I__7970 (
            .O(N__38390),
            .I(N__38385));
    InMux I__7969 (
            .O(N__38389),
            .I(N__38382));
    InMux I__7968 (
            .O(N__38388),
            .I(N__38377));
    InMux I__7967 (
            .O(N__38385),
            .I(N__38377));
    LocalMux I__7966 (
            .O(N__38382),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__7965 (
            .O(N__38377),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    CascadeMux I__7964 (
            .O(N__38372),
            .I(N__38369));
    InMux I__7963 (
            .O(N__38369),
            .I(N__38366));
    LocalMux I__7962 (
            .O(N__38366),
            .I(N__38363));
    Span4Mux_h I__7961 (
            .O(N__38363),
            .I(N__38360));
    Odrv4 I__7960 (
            .O(N__38360),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt28 ));
    InMux I__7959 (
            .O(N__38357),
            .I(N__38354));
    LocalMux I__7958 (
            .O(N__38354),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__7957 (
            .O(N__38351),
            .I(N__38348));
    InMux I__7956 (
            .O(N__38348),
            .I(N__38345));
    LocalMux I__7955 (
            .O(N__38345),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    InMux I__7954 (
            .O(N__38342),
            .I(N__38338));
    InMux I__7953 (
            .O(N__38341),
            .I(N__38335));
    LocalMux I__7952 (
            .O(N__38338),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    LocalMux I__7951 (
            .O(N__38335),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    InMux I__7950 (
            .O(N__38330),
            .I(N__38327));
    LocalMux I__7949 (
            .O(N__38327),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    InMux I__7948 (
            .O(N__38324),
            .I(N__38321));
    LocalMux I__7947 (
            .O(N__38321),
            .I(N__38318));
    Span4Mux_h I__7946 (
            .O(N__38318),
            .I(N__38315));
    Odrv4 I__7945 (
            .O(N__38315),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__7944 (
            .O(N__38312),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ));
    InMux I__7943 (
            .O(N__38309),
            .I(N__38306));
    LocalMux I__7942 (
            .O(N__38306),
            .I(N__38303));
    Odrv12 I__7941 (
            .O(N__38303),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    InMux I__7940 (
            .O(N__38300),
            .I(N__38296));
    InMux I__7939 (
            .O(N__38299),
            .I(N__38293));
    LocalMux I__7938 (
            .O(N__38296),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    LocalMux I__7937 (
            .O(N__38293),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    InMux I__7936 (
            .O(N__38288),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__7935 (
            .O(N__38285),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__7934 (
            .O(N__38282),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__7933 (
            .O(N__38279),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__7932 (
            .O(N__38276),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__7931 (
            .O(N__38273),
            .I(N__38270));
    LocalMux I__7930 (
            .O(N__38270),
            .I(N__38267));
    Span4Mux_v I__7929 (
            .O(N__38267),
            .I(N__38264));
    Odrv4 I__7928 (
            .O(N__38264),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    InMux I__7927 (
            .O(N__38261),
            .I(N__38256));
    InMux I__7926 (
            .O(N__38260),
            .I(N__38251));
    InMux I__7925 (
            .O(N__38259),
            .I(N__38251));
    LocalMux I__7924 (
            .O(N__38256),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__7923 (
            .O(N__38251),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__7922 (
            .O(N__38246),
            .I(N__38243));
    InMux I__7921 (
            .O(N__38243),
            .I(N__38236));
    InMux I__7920 (
            .O(N__38242),
            .I(N__38236));
    InMux I__7919 (
            .O(N__38241),
            .I(N__38233));
    LocalMux I__7918 (
            .O(N__38236),
            .I(N__38230));
    LocalMux I__7917 (
            .O(N__38233),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__7916 (
            .O(N__38230),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__7915 (
            .O(N__38225),
            .I(N__38222));
    InMux I__7914 (
            .O(N__38222),
            .I(N__38219));
    LocalMux I__7913 (
            .O(N__38219),
            .I(N__38216));
    Span4Mux_v I__7912 (
            .O(N__38216),
            .I(N__38213));
    Odrv4 I__7911 (
            .O(N__38213),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    InMux I__7910 (
            .O(N__38210),
            .I(N__38204));
    InMux I__7909 (
            .O(N__38209),
            .I(N__38204));
    LocalMux I__7908 (
            .O(N__38204),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__7907 (
            .O(N__38201),
            .I(N__38198));
    InMux I__7906 (
            .O(N__38198),
            .I(N__38192));
    InMux I__7905 (
            .O(N__38197),
            .I(N__38192));
    LocalMux I__7904 (
            .O(N__38192),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    InMux I__7903 (
            .O(N__38189),
            .I(bfn_15_19_0_));
    InMux I__7902 (
            .O(N__38186),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__7901 (
            .O(N__38183),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__7900 (
            .O(N__38180),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__7899 (
            .O(N__38177),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__7898 (
            .O(N__38174),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__7897 (
            .O(N__38171),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__7896 (
            .O(N__38168),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__7895 (
            .O(N__38165),
            .I(bfn_15_20_0_));
    InMux I__7894 (
            .O(N__38162),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__7893 (
            .O(N__38159),
            .I(bfn_15_18_0_));
    InMux I__7892 (
            .O(N__38156),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__7891 (
            .O(N__38153),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__7890 (
            .O(N__38150),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__7889 (
            .O(N__38147),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__7888 (
            .O(N__38144),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__7887 (
            .O(N__38141),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__7886 (
            .O(N__38138),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__7885 (
            .O(N__38135),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__7884 (
            .O(N__38132),
            .I(N__38108));
    InMux I__7883 (
            .O(N__38131),
            .I(N__38108));
    InMux I__7882 (
            .O(N__38130),
            .I(N__38108));
    InMux I__7881 (
            .O(N__38129),
            .I(N__38108));
    InMux I__7880 (
            .O(N__38128),
            .I(N__38099));
    InMux I__7879 (
            .O(N__38127),
            .I(N__38099));
    InMux I__7878 (
            .O(N__38126),
            .I(N__38099));
    InMux I__7877 (
            .O(N__38125),
            .I(N__38099));
    InMux I__7876 (
            .O(N__38124),
            .I(N__38076));
    InMux I__7875 (
            .O(N__38123),
            .I(N__38076));
    InMux I__7874 (
            .O(N__38122),
            .I(N__38076));
    InMux I__7873 (
            .O(N__38121),
            .I(N__38076));
    InMux I__7872 (
            .O(N__38120),
            .I(N__38067));
    InMux I__7871 (
            .O(N__38119),
            .I(N__38067));
    InMux I__7870 (
            .O(N__38118),
            .I(N__38067));
    InMux I__7869 (
            .O(N__38117),
            .I(N__38067));
    LocalMux I__7868 (
            .O(N__38108),
            .I(N__38062));
    LocalMux I__7867 (
            .O(N__38099),
            .I(N__38062));
    InMux I__7866 (
            .O(N__38098),
            .I(N__38053));
    InMux I__7865 (
            .O(N__38097),
            .I(N__38053));
    InMux I__7864 (
            .O(N__38096),
            .I(N__38053));
    InMux I__7863 (
            .O(N__38095),
            .I(N__38053));
    InMux I__7862 (
            .O(N__38094),
            .I(N__38048));
    InMux I__7861 (
            .O(N__38093),
            .I(N__38048));
    InMux I__7860 (
            .O(N__38092),
            .I(N__38039));
    InMux I__7859 (
            .O(N__38091),
            .I(N__38039));
    InMux I__7858 (
            .O(N__38090),
            .I(N__38039));
    InMux I__7857 (
            .O(N__38089),
            .I(N__38039));
    InMux I__7856 (
            .O(N__38088),
            .I(N__38030));
    InMux I__7855 (
            .O(N__38087),
            .I(N__38030));
    InMux I__7854 (
            .O(N__38086),
            .I(N__38030));
    InMux I__7853 (
            .O(N__38085),
            .I(N__38030));
    LocalMux I__7852 (
            .O(N__38076),
            .I(N__38025));
    LocalMux I__7851 (
            .O(N__38067),
            .I(N__38025));
    Span4Mux_v I__7850 (
            .O(N__38062),
            .I(N__38014));
    LocalMux I__7849 (
            .O(N__38053),
            .I(N__38014));
    LocalMux I__7848 (
            .O(N__38048),
            .I(N__38014));
    LocalMux I__7847 (
            .O(N__38039),
            .I(N__38014));
    LocalMux I__7846 (
            .O(N__38030),
            .I(N__38014));
    Span4Mux_v I__7845 (
            .O(N__38025),
            .I(N__38009));
    Span4Mux_v I__7844 (
            .O(N__38014),
            .I(N__38009));
    Odrv4 I__7843 (
            .O(N__38009),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__7842 (
            .O(N__38006),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CEMux I__7841 (
            .O(N__38003),
            .I(N__37998));
    CEMux I__7840 (
            .O(N__38002),
            .I(N__37995));
    CEMux I__7839 (
            .O(N__38001),
            .I(N__37992));
    LocalMux I__7838 (
            .O(N__37998),
            .I(N__37988));
    LocalMux I__7837 (
            .O(N__37995),
            .I(N__37983));
    LocalMux I__7836 (
            .O(N__37992),
            .I(N__37983));
    CEMux I__7835 (
            .O(N__37991),
            .I(N__37980));
    Span4Mux_v I__7834 (
            .O(N__37988),
            .I(N__37973));
    Span4Mux_v I__7833 (
            .O(N__37983),
            .I(N__37973));
    LocalMux I__7832 (
            .O(N__37980),
            .I(N__37973));
    Span4Mux_v I__7831 (
            .O(N__37973),
            .I(N__37970));
    Span4Mux_h I__7830 (
            .O(N__37970),
            .I(N__37967));
    Odrv4 I__7829 (
            .O(N__37967),
            .I(\current_shift_inst.timer_s1.N_168_i ));
    InMux I__7828 (
            .O(N__37964),
            .I(bfn_15_17_0_));
    InMux I__7827 (
            .O(N__37961),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__7826 (
            .O(N__37958),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__7825 (
            .O(N__37955),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__7824 (
            .O(N__37952),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__7823 (
            .O(N__37949),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__7822 (
            .O(N__37946),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__7821 (
            .O(N__37943),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__7820 (
            .O(N__37940),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__7819 (
            .O(N__37937),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__7818 (
            .O(N__37934),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__7817 (
            .O(N__37931),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__7816 (
            .O(N__37928),
            .I(bfn_15_16_0_));
    InMux I__7815 (
            .O(N__37925),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__7814 (
            .O(N__37922),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__7813 (
            .O(N__37919),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__7812 (
            .O(N__37916),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__7811 (
            .O(N__37913),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__7810 (
            .O(N__37910),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    InMux I__7809 (
            .O(N__37907),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__7808 (
            .O(N__37904),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__7807 (
            .O(N__37901),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    InMux I__7806 (
            .O(N__37898),
            .I(bfn_15_15_0_));
    InMux I__7805 (
            .O(N__37895),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__7804 (
            .O(N__37892),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__7803 (
            .O(N__37889),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__7802 (
            .O(N__37886),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__7801 (
            .O(N__37883),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__7800 (
            .O(N__37880),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    InMux I__7799 (
            .O(N__37877),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__7798 (
            .O(N__37874),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__7797 (
            .O(N__37871),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    InMux I__7796 (
            .O(N__37868),
            .I(bfn_15_14_0_));
    InMux I__7795 (
            .O(N__37865),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__7794 (
            .O(N__37862),
            .I(N__37859));
    InMux I__7793 (
            .O(N__37859),
            .I(N__37856));
    LocalMux I__7792 (
            .O(N__37856),
            .I(N__37853));
    Odrv4 I__7791 (
            .O(N__37853),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    CascadeMux I__7790 (
            .O(N__37850),
            .I(N__37847));
    InMux I__7789 (
            .O(N__37847),
            .I(N__37844));
    LocalMux I__7788 (
            .O(N__37844),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__7787 (
            .O(N__37841),
            .I(N__37838));
    LocalMux I__7786 (
            .O(N__37838),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__7785 (
            .O(N__37835),
            .I(N__37832));
    LocalMux I__7784 (
            .O(N__37832),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    CascadeMux I__7783 (
            .O(N__37829),
            .I(N__37826));
    InMux I__7782 (
            .O(N__37826),
            .I(N__37823));
    LocalMux I__7781 (
            .O(N__37823),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    CascadeMux I__7780 (
            .O(N__37820),
            .I(N__37817));
    InMux I__7779 (
            .O(N__37817),
            .I(N__37814));
    LocalMux I__7778 (
            .O(N__37814),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    CascadeMux I__7777 (
            .O(N__37811),
            .I(N__37808));
    InMux I__7776 (
            .O(N__37808),
            .I(N__37805));
    LocalMux I__7775 (
            .O(N__37805),
            .I(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ));
    InMux I__7774 (
            .O(N__37802),
            .I(N__37799));
    LocalMux I__7773 (
            .O(N__37799),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__7772 (
            .O(N__37796),
            .I(bfn_15_13_0_));
    CascadeMux I__7771 (
            .O(N__37793),
            .I(N__37790));
    InMux I__7770 (
            .O(N__37790),
            .I(N__37787));
    LocalMux I__7769 (
            .O(N__37787),
            .I(N__37784));
    Odrv4 I__7768 (
            .O(N__37784),
            .I(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ));
    InMux I__7767 (
            .O(N__37781),
            .I(N__37778));
    LocalMux I__7766 (
            .O(N__37778),
            .I(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ));
    InMux I__7765 (
            .O(N__37775),
            .I(N__37772));
    LocalMux I__7764 (
            .O(N__37772),
            .I(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ));
    InMux I__7763 (
            .O(N__37769),
            .I(N__37766));
    LocalMux I__7762 (
            .O(N__37766),
            .I(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ));
    CascadeMux I__7761 (
            .O(N__37763),
            .I(N__37760));
    InMux I__7760 (
            .O(N__37760),
            .I(N__37757));
    LocalMux I__7759 (
            .O(N__37757),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__7758 (
            .O(N__37754),
            .I(N__37751));
    LocalMux I__7757 (
            .O(N__37751),
            .I(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ));
    CascadeMux I__7756 (
            .O(N__37748),
            .I(N__37745));
    InMux I__7755 (
            .O(N__37745),
            .I(N__37742));
    LocalMux I__7754 (
            .O(N__37742),
            .I(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ));
    CascadeMux I__7753 (
            .O(N__37739),
            .I(N__37736));
    InMux I__7752 (
            .O(N__37736),
            .I(N__37733));
    LocalMux I__7751 (
            .O(N__37733),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__7750 (
            .O(N__37730),
            .I(N__37727));
    LocalMux I__7749 (
            .O(N__37727),
            .I(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ));
    CascadeMux I__7748 (
            .O(N__37724),
            .I(N__37721));
    InMux I__7747 (
            .O(N__37721),
            .I(N__37718));
    LocalMux I__7746 (
            .O(N__37718),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    CascadeMux I__7745 (
            .O(N__37715),
            .I(N__37712));
    InMux I__7744 (
            .O(N__37712),
            .I(N__37709));
    LocalMux I__7743 (
            .O(N__37709),
            .I(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ));
    CascadeMux I__7742 (
            .O(N__37706),
            .I(N__37703));
    InMux I__7741 (
            .O(N__37703),
            .I(N__37700));
    LocalMux I__7740 (
            .O(N__37700),
            .I(N__37697));
    Odrv4 I__7739 (
            .O(N__37697),
            .I(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ));
    CascadeMux I__7738 (
            .O(N__37694),
            .I(N__37691));
    InMux I__7737 (
            .O(N__37691),
            .I(N__37688));
    LocalMux I__7736 (
            .O(N__37688),
            .I(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ));
    CascadeMux I__7735 (
            .O(N__37685),
            .I(N__37682));
    InMux I__7734 (
            .O(N__37682),
            .I(N__37679));
    LocalMux I__7733 (
            .O(N__37679),
            .I(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ));
    InMux I__7732 (
            .O(N__37676),
            .I(N__37673));
    LocalMux I__7731 (
            .O(N__37673),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__7730 (
            .O(N__37670),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__7729 (
            .O(N__37667),
            .I(N__37661));
    InMux I__7728 (
            .O(N__37666),
            .I(N__37658));
    InMux I__7727 (
            .O(N__37665),
            .I(N__37653));
    InMux I__7726 (
            .O(N__37664),
            .I(N__37653));
    LocalMux I__7725 (
            .O(N__37661),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__7724 (
            .O(N__37658),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__7723 (
            .O(N__37653),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__7722 (
            .O(N__37646),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    CascadeMux I__7721 (
            .O(N__37643),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    CascadeMux I__7720 (
            .O(N__37640),
            .I(N__37637));
    InMux I__7719 (
            .O(N__37637),
            .I(N__37633));
    InMux I__7718 (
            .O(N__37636),
            .I(N__37630));
    LocalMux I__7717 (
            .O(N__37633),
            .I(N__37627));
    LocalMux I__7716 (
            .O(N__37630),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv4 I__7715 (
            .O(N__37627),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    InMux I__7714 (
            .O(N__37622),
            .I(N__37619));
    LocalMux I__7713 (
            .O(N__37619),
            .I(N__37616));
    Span4Mux_v I__7712 (
            .O(N__37616),
            .I(N__37612));
    InMux I__7711 (
            .O(N__37615),
            .I(N__37609));
    Odrv4 I__7710 (
            .O(N__37612),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    LocalMux I__7709 (
            .O(N__37609),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    InMux I__7708 (
            .O(N__37604),
            .I(N__37601));
    LocalMux I__7707 (
            .O(N__37601),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CascadeMux I__7706 (
            .O(N__37598),
            .I(N__37595));
    InMux I__7705 (
            .O(N__37595),
            .I(N__37592));
    LocalMux I__7704 (
            .O(N__37592),
            .I(N__37587));
    CascadeMux I__7703 (
            .O(N__37591),
            .I(N__37584));
    InMux I__7702 (
            .O(N__37590),
            .I(N__37580));
    Span4Mux_v I__7701 (
            .O(N__37587),
            .I(N__37577));
    InMux I__7700 (
            .O(N__37584),
            .I(N__37574));
    InMux I__7699 (
            .O(N__37583),
            .I(N__37571));
    LocalMux I__7698 (
            .O(N__37580),
            .I(N__37568));
    Odrv4 I__7697 (
            .O(N__37577),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__7696 (
            .O(N__37574),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__7695 (
            .O(N__37571),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv12 I__7694 (
            .O(N__37568),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__7693 (
            .O(N__37559),
            .I(N__37556));
    InMux I__7692 (
            .O(N__37556),
            .I(N__37553));
    LocalMux I__7691 (
            .O(N__37553),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__7690 (
            .O(N__37550),
            .I(N__37547));
    LocalMux I__7689 (
            .O(N__37547),
            .I(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ));
    InMux I__7688 (
            .O(N__37544),
            .I(N__37541));
    LocalMux I__7687 (
            .O(N__37541),
            .I(N__37538));
    Span4Mux_v I__7686 (
            .O(N__37538),
            .I(N__37535));
    Odrv4 I__7685 (
            .O(N__37535),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    CascadeMux I__7684 (
            .O(N__37532),
            .I(N__37529));
    InMux I__7683 (
            .O(N__37529),
            .I(N__37526));
    LocalMux I__7682 (
            .O(N__37526),
            .I(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ));
    InMux I__7681 (
            .O(N__37523),
            .I(N__37520));
    LocalMux I__7680 (
            .O(N__37520),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    InMux I__7679 (
            .O(N__37517),
            .I(N__37514));
    LocalMux I__7678 (
            .O(N__37514),
            .I(N__37511));
    Odrv4 I__7677 (
            .O(N__37511),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    CascadeMux I__7676 (
            .O(N__37508),
            .I(N__37505));
    InMux I__7675 (
            .O(N__37505),
            .I(N__37502));
    LocalMux I__7674 (
            .O(N__37502),
            .I(N__37499));
    Odrv4 I__7673 (
            .O(N__37499),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    CascadeMux I__7672 (
            .O(N__37496),
            .I(N__37493));
    InMux I__7671 (
            .O(N__37493),
            .I(N__37490));
    LocalMux I__7670 (
            .O(N__37490),
            .I(N__37487));
    Odrv4 I__7669 (
            .O(N__37487),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    CascadeMux I__7668 (
            .O(N__37484),
            .I(N__37481));
    InMux I__7667 (
            .O(N__37481),
            .I(N__37478));
    LocalMux I__7666 (
            .O(N__37478),
            .I(N__37475));
    Span4Mux_h I__7665 (
            .O(N__37475),
            .I(N__37472));
    Odrv4 I__7664 (
            .O(N__37472),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__7663 (
            .O(N__37469),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__7662 (
            .O(N__37466),
            .I(N__37463));
    InMux I__7661 (
            .O(N__37463),
            .I(N__37460));
    LocalMux I__7660 (
            .O(N__37460),
            .I(N__37457));
    Odrv12 I__7659 (
            .O(N__37457),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    CascadeMux I__7658 (
            .O(N__37454),
            .I(N__37451));
    InMux I__7657 (
            .O(N__37451),
            .I(N__37448));
    LocalMux I__7656 (
            .O(N__37448),
            .I(N__37445));
    Span4Mux_h I__7655 (
            .O(N__37445),
            .I(N__37442));
    Span4Mux_v I__7654 (
            .O(N__37442),
            .I(N__37439));
    Odrv4 I__7653 (
            .O(N__37439),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ));
    IoInMux I__7652 (
            .O(N__37436),
            .I(N__37410));
    InMux I__7651 (
            .O(N__37435),
            .I(N__37393));
    InMux I__7650 (
            .O(N__37434),
            .I(N__37393));
    InMux I__7649 (
            .O(N__37433),
            .I(N__37393));
    InMux I__7648 (
            .O(N__37432),
            .I(N__37393));
    InMux I__7647 (
            .O(N__37431),
            .I(N__37384));
    InMux I__7646 (
            .O(N__37430),
            .I(N__37384));
    InMux I__7645 (
            .O(N__37429),
            .I(N__37384));
    InMux I__7644 (
            .O(N__37428),
            .I(N__37384));
    InMux I__7643 (
            .O(N__37427),
            .I(N__37377));
    InMux I__7642 (
            .O(N__37426),
            .I(N__37377));
    InMux I__7641 (
            .O(N__37425),
            .I(N__37377));
    InMux I__7640 (
            .O(N__37424),
            .I(N__37368));
    InMux I__7639 (
            .O(N__37423),
            .I(N__37368));
    InMux I__7638 (
            .O(N__37422),
            .I(N__37368));
    InMux I__7637 (
            .O(N__37421),
            .I(N__37368));
    InMux I__7636 (
            .O(N__37420),
            .I(N__37359));
    InMux I__7635 (
            .O(N__37419),
            .I(N__37359));
    InMux I__7634 (
            .O(N__37418),
            .I(N__37359));
    InMux I__7633 (
            .O(N__37417),
            .I(N__37359));
    InMux I__7632 (
            .O(N__37416),
            .I(N__37350));
    InMux I__7631 (
            .O(N__37415),
            .I(N__37350));
    InMux I__7630 (
            .O(N__37414),
            .I(N__37350));
    InMux I__7629 (
            .O(N__37413),
            .I(N__37350));
    LocalMux I__7628 (
            .O(N__37410),
            .I(N__37347));
    InMux I__7627 (
            .O(N__37409),
            .I(N__37344));
    InMux I__7626 (
            .O(N__37408),
            .I(N__37337));
    InMux I__7625 (
            .O(N__37407),
            .I(N__37337));
    InMux I__7624 (
            .O(N__37406),
            .I(N__37337));
    InMux I__7623 (
            .O(N__37405),
            .I(N__37328));
    InMux I__7622 (
            .O(N__37404),
            .I(N__37328));
    InMux I__7621 (
            .O(N__37403),
            .I(N__37328));
    InMux I__7620 (
            .O(N__37402),
            .I(N__37328));
    LocalMux I__7619 (
            .O(N__37393),
            .I(N__37323));
    LocalMux I__7618 (
            .O(N__37384),
            .I(N__37323));
    LocalMux I__7617 (
            .O(N__37377),
            .I(N__37314));
    LocalMux I__7616 (
            .O(N__37368),
            .I(N__37314));
    LocalMux I__7615 (
            .O(N__37359),
            .I(N__37314));
    LocalMux I__7614 (
            .O(N__37350),
            .I(N__37314));
    Span4Mux_s1_v I__7613 (
            .O(N__37347),
            .I(N__37311));
    LocalMux I__7612 (
            .O(N__37344),
            .I(N__37308));
    LocalMux I__7611 (
            .O(N__37337),
            .I(N__37299));
    LocalMux I__7610 (
            .O(N__37328),
            .I(N__37299));
    Span4Mux_v I__7609 (
            .O(N__37323),
            .I(N__37299));
    Span4Mux_v I__7608 (
            .O(N__37314),
            .I(N__37299));
    Span4Mux_h I__7607 (
            .O(N__37311),
            .I(N__37296));
    Span4Mux_v I__7606 (
            .O(N__37308),
            .I(N__37289));
    Span4Mux_v I__7605 (
            .O(N__37299),
            .I(N__37289));
    Span4Mux_v I__7604 (
            .O(N__37296),
            .I(N__37289));
    Odrv4 I__7603 (
            .O(N__37289),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__7602 (
            .O(N__37286),
            .I(N__37280));
    InMux I__7601 (
            .O(N__37285),
            .I(N__37280));
    LocalMux I__7600 (
            .O(N__37280),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__7599 (
            .O(N__37277),
            .I(N__37274));
    InMux I__7598 (
            .O(N__37274),
            .I(N__37270));
    InMux I__7597 (
            .O(N__37273),
            .I(N__37264));
    LocalMux I__7596 (
            .O(N__37270),
            .I(N__37261));
    InMux I__7595 (
            .O(N__37269),
            .I(N__37254));
    InMux I__7594 (
            .O(N__37268),
            .I(N__37254));
    InMux I__7593 (
            .O(N__37267),
            .I(N__37254));
    LocalMux I__7592 (
            .O(N__37264),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__7591 (
            .O(N__37261),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    LocalMux I__7590 (
            .O(N__37254),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__7589 (
            .O(N__37247),
            .I(N__37244));
    LocalMux I__7588 (
            .O(N__37244),
            .I(N__37239));
    InMux I__7587 (
            .O(N__37243),
            .I(N__37236));
    CascadeMux I__7586 (
            .O(N__37242),
            .I(N__37233));
    Span4Mux_v I__7585 (
            .O(N__37239),
            .I(N__37228));
    LocalMux I__7584 (
            .O(N__37236),
            .I(N__37228));
    InMux I__7583 (
            .O(N__37233),
            .I(N__37225));
    Span4Mux_v I__7582 (
            .O(N__37228),
            .I(N__37222));
    LocalMux I__7581 (
            .O(N__37225),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__7580 (
            .O(N__37222),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__7579 (
            .O(N__37217),
            .I(N__37214));
    InMux I__7578 (
            .O(N__37214),
            .I(N__37211));
    LocalMux I__7577 (
            .O(N__37211),
            .I(N__37208));
    Odrv4 I__7576 (
            .O(N__37208),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    CascadeMux I__7575 (
            .O(N__37205),
            .I(N__37202));
    InMux I__7574 (
            .O(N__37202),
            .I(N__37199));
    LocalMux I__7573 (
            .O(N__37199),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    CascadeMux I__7572 (
            .O(N__37196),
            .I(N__37193));
    InMux I__7571 (
            .O(N__37193),
            .I(N__37190));
    LocalMux I__7570 (
            .O(N__37190),
            .I(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ));
    CascadeMux I__7569 (
            .O(N__37187),
            .I(N__37184));
    InMux I__7568 (
            .O(N__37184),
            .I(N__37181));
    LocalMux I__7567 (
            .O(N__37181),
            .I(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ));
    CascadeMux I__7566 (
            .O(N__37178),
            .I(N__37175));
    InMux I__7565 (
            .O(N__37175),
            .I(N__37172));
    LocalMux I__7564 (
            .O(N__37172),
            .I(N__37169));
    Odrv4 I__7563 (
            .O(N__37169),
            .I(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ));
    InMux I__7562 (
            .O(N__37166),
            .I(N__37163));
    LocalMux I__7561 (
            .O(N__37163),
            .I(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ));
    InMux I__7560 (
            .O(N__37160),
            .I(N__37157));
    LocalMux I__7559 (
            .O(N__37157),
            .I(N__37154));
    Span4Mux_v I__7558 (
            .O(N__37154),
            .I(N__37151));
    Odrv4 I__7557 (
            .O(N__37151),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ));
    CascadeMux I__7556 (
            .O(N__37148),
            .I(N__37145));
    InMux I__7555 (
            .O(N__37145),
            .I(N__37142));
    LocalMux I__7554 (
            .O(N__37142),
            .I(N__37139));
    Span4Mux_v I__7553 (
            .O(N__37139),
            .I(N__37136));
    Odrv4 I__7552 (
            .O(N__37136),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt20 ));
    InMux I__7551 (
            .O(N__37133),
            .I(N__37130));
    LocalMux I__7550 (
            .O(N__37130),
            .I(N__37127));
    Span4Mux_v I__7549 (
            .O(N__37127),
            .I(N__37124));
    Odrv4 I__7548 (
            .O(N__37124),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ));
    CascadeMux I__7547 (
            .O(N__37121),
            .I(N__37118));
    InMux I__7546 (
            .O(N__37118),
            .I(N__37115));
    LocalMux I__7545 (
            .O(N__37115),
            .I(N__37112));
    Span4Mux_h I__7544 (
            .O(N__37112),
            .I(N__37109));
    Span4Mux_v I__7543 (
            .O(N__37109),
            .I(N__37106));
    Odrv4 I__7542 (
            .O(N__37106),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt22 ));
    InMux I__7541 (
            .O(N__37103),
            .I(N__37100));
    LocalMux I__7540 (
            .O(N__37100),
            .I(N__37097));
    Odrv12 I__7539 (
            .O(N__37097),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt24 ));
    CascadeMux I__7538 (
            .O(N__37094),
            .I(N__37091));
    InMux I__7537 (
            .O(N__37091),
            .I(N__37088));
    LocalMux I__7536 (
            .O(N__37088),
            .I(N__37085));
    Odrv12 I__7535 (
            .O(N__37085),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ));
    InMux I__7534 (
            .O(N__37082),
            .I(N__37079));
    LocalMux I__7533 (
            .O(N__37079),
            .I(N__37076));
    Odrv4 I__7532 (
            .O(N__37076),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ));
    InMux I__7531 (
            .O(N__37073),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ));
    InMux I__7530 (
            .O(N__37070),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    InMux I__7529 (
            .O(N__37067),
            .I(N__37063));
    InMux I__7528 (
            .O(N__37066),
            .I(N__37060));
    LocalMux I__7527 (
            .O(N__37063),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    LocalMux I__7526 (
            .O(N__37060),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__7525 (
            .O(N__37055),
            .I(N__37052));
    LocalMux I__7524 (
            .O(N__37052),
            .I(N__37045));
    InMux I__7523 (
            .O(N__37051),
            .I(N__37042));
    InMux I__7522 (
            .O(N__37050),
            .I(N__37039));
    InMux I__7521 (
            .O(N__37049),
            .I(N__37036));
    InMux I__7520 (
            .O(N__37048),
            .I(N__37033));
    Span4Mux_h I__7519 (
            .O(N__37045),
            .I(N__37030));
    LocalMux I__7518 (
            .O(N__37042),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__7517 (
            .O(N__37039),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__7516 (
            .O(N__37036),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__7515 (
            .O(N__37033),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__7514 (
            .O(N__37030),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    CascadeMux I__7513 (
            .O(N__37019),
            .I(N__37016));
    InMux I__7512 (
            .O(N__37016),
            .I(N__37013));
    LocalMux I__7511 (
            .O(N__37013),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df30 ));
    InMux I__7510 (
            .O(N__37010),
            .I(N__37007));
    LocalMux I__7509 (
            .O(N__37007),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__7508 (
            .O(N__37004),
            .I(N__37000));
    InMux I__7507 (
            .O(N__37003),
            .I(N__36997));
    LocalMux I__7506 (
            .O(N__37000),
            .I(N__36994));
    LocalMux I__7505 (
            .O(N__36997),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv12 I__7504 (
            .O(N__36994),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__7503 (
            .O(N__36989),
            .I(N__36986));
    LocalMux I__7502 (
            .O(N__36986),
            .I(N__36983));
    Span4Mux_v I__7501 (
            .O(N__36983),
            .I(N__36980));
    Odrv4 I__7500 (
            .O(N__36980),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__7499 (
            .O(N__36977),
            .I(N__36974));
    InMux I__7498 (
            .O(N__36974),
            .I(N__36971));
    LocalMux I__7497 (
            .O(N__36971),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__7496 (
            .O(N__36968),
            .I(N__36965));
    LocalMux I__7495 (
            .O(N__36965),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    InMux I__7494 (
            .O(N__36962),
            .I(N__36958));
    InMux I__7493 (
            .O(N__36961),
            .I(N__36955));
    LocalMux I__7492 (
            .O(N__36958),
            .I(N__36952));
    LocalMux I__7491 (
            .O(N__36955),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv12 I__7490 (
            .O(N__36952),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__7489 (
            .O(N__36947),
            .I(N__36944));
    InMux I__7488 (
            .O(N__36944),
            .I(N__36941));
    LocalMux I__7487 (
            .O(N__36941),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__7486 (
            .O(N__36938),
            .I(N__36935));
    InMux I__7485 (
            .O(N__36935),
            .I(N__36932));
    LocalMux I__7484 (
            .O(N__36932),
            .I(N__36929));
    Odrv12 I__7483 (
            .O(N__36929),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__7482 (
            .O(N__36926),
            .I(N__36922));
    InMux I__7481 (
            .O(N__36925),
            .I(N__36919));
    LocalMux I__7480 (
            .O(N__36922),
            .I(N__36916));
    LocalMux I__7479 (
            .O(N__36919),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv12 I__7478 (
            .O(N__36916),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__7477 (
            .O(N__36911),
            .I(N__36908));
    LocalMux I__7476 (
            .O(N__36908),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__7475 (
            .O(N__36905),
            .I(N__36902));
    InMux I__7474 (
            .O(N__36902),
            .I(N__36899));
    LocalMux I__7473 (
            .O(N__36899),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__7472 (
            .O(N__36896),
            .I(N__36893));
    LocalMux I__7471 (
            .O(N__36893),
            .I(N__36889));
    InMux I__7470 (
            .O(N__36892),
            .I(N__36886));
    Span4Mux_v I__7469 (
            .O(N__36889),
            .I(N__36883));
    LocalMux I__7468 (
            .O(N__36886),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__7467 (
            .O(N__36883),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__7466 (
            .O(N__36878),
            .I(N__36875));
    LocalMux I__7465 (
            .O(N__36875),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__7464 (
            .O(N__36872),
            .I(N__36869));
    LocalMux I__7463 (
            .O(N__36869),
            .I(N__36866));
    Span4Mux_v I__7462 (
            .O(N__36866),
            .I(N__36863));
    Span4Mux_v I__7461 (
            .O(N__36863),
            .I(N__36860));
    Odrv4 I__7460 (
            .O(N__36860),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    InMux I__7459 (
            .O(N__36857),
            .I(N__36853));
    InMux I__7458 (
            .O(N__36856),
            .I(N__36850));
    LocalMux I__7457 (
            .O(N__36853),
            .I(N__36847));
    LocalMux I__7456 (
            .O(N__36850),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv12 I__7455 (
            .O(N__36847),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__7454 (
            .O(N__36842),
            .I(N__36839));
    InMux I__7453 (
            .O(N__36839),
            .I(N__36836));
    LocalMux I__7452 (
            .O(N__36836),
            .I(N__36833));
    Odrv4 I__7451 (
            .O(N__36833),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__7450 (
            .O(N__36830),
            .I(N__36826));
    InMux I__7449 (
            .O(N__36829),
            .I(N__36823));
    LocalMux I__7448 (
            .O(N__36826),
            .I(N__36820));
    LocalMux I__7447 (
            .O(N__36823),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv12 I__7446 (
            .O(N__36820),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__7445 (
            .O(N__36815),
            .I(N__36812));
    LocalMux I__7444 (
            .O(N__36812),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__7443 (
            .O(N__36809),
            .I(N__36806));
    LocalMux I__7442 (
            .O(N__36806),
            .I(N__36802));
    InMux I__7441 (
            .O(N__36805),
            .I(N__36799));
    Span4Mux_v I__7440 (
            .O(N__36802),
            .I(N__36796));
    LocalMux I__7439 (
            .O(N__36799),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__7438 (
            .O(N__36796),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__7437 (
            .O(N__36791),
            .I(N__36788));
    LocalMux I__7436 (
            .O(N__36788),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__7435 (
            .O(N__36785),
            .I(N__36782));
    LocalMux I__7434 (
            .O(N__36782),
            .I(N__36778));
    InMux I__7433 (
            .O(N__36781),
            .I(N__36775));
    Span4Mux_v I__7432 (
            .O(N__36778),
            .I(N__36772));
    LocalMux I__7431 (
            .O(N__36775),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__7430 (
            .O(N__36772),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__7429 (
            .O(N__36767),
            .I(N__36764));
    InMux I__7428 (
            .O(N__36764),
            .I(N__36761));
    LocalMux I__7427 (
            .O(N__36761),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__7426 (
            .O(N__36758),
            .I(N__36755));
    LocalMux I__7425 (
            .O(N__36755),
            .I(N__36751));
    InMux I__7424 (
            .O(N__36754),
            .I(N__36748));
    Span4Mux_v I__7423 (
            .O(N__36751),
            .I(N__36745));
    LocalMux I__7422 (
            .O(N__36748),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__7421 (
            .O(N__36745),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__7420 (
            .O(N__36740),
            .I(N__36737));
    InMux I__7419 (
            .O(N__36737),
            .I(N__36734));
    LocalMux I__7418 (
            .O(N__36734),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__7417 (
            .O(N__36731),
            .I(N__36727));
    InMux I__7416 (
            .O(N__36730),
            .I(N__36724));
    LocalMux I__7415 (
            .O(N__36727),
            .I(N__36721));
    LocalMux I__7414 (
            .O(N__36724),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv12 I__7413 (
            .O(N__36721),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__7412 (
            .O(N__36716),
            .I(N__36713));
    InMux I__7411 (
            .O(N__36713),
            .I(N__36710));
    LocalMux I__7410 (
            .O(N__36710),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__7409 (
            .O(N__36707),
            .I(N__36704));
    LocalMux I__7408 (
            .O(N__36704),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__7407 (
            .O(N__36701),
            .I(N__36697));
    InMux I__7406 (
            .O(N__36700),
            .I(N__36694));
    LocalMux I__7405 (
            .O(N__36697),
            .I(N__36691));
    LocalMux I__7404 (
            .O(N__36694),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv12 I__7403 (
            .O(N__36691),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__7402 (
            .O(N__36686),
            .I(N__36683));
    InMux I__7401 (
            .O(N__36683),
            .I(N__36680));
    LocalMux I__7400 (
            .O(N__36680),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__7399 (
            .O(N__36677),
            .I(N__36674));
    LocalMux I__7398 (
            .O(N__36674),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    InMux I__7397 (
            .O(N__36671),
            .I(N__36667));
    InMux I__7396 (
            .O(N__36670),
            .I(N__36664));
    LocalMux I__7395 (
            .O(N__36667),
            .I(N__36661));
    LocalMux I__7394 (
            .O(N__36664),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv12 I__7393 (
            .O(N__36661),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__7392 (
            .O(N__36656),
            .I(N__36653));
    InMux I__7391 (
            .O(N__36653),
            .I(N__36650));
    LocalMux I__7390 (
            .O(N__36650),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__7389 (
            .O(N__36647),
            .I(N__36644));
    LocalMux I__7388 (
            .O(N__36644),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    InMux I__7387 (
            .O(N__36641),
            .I(N__36637));
    InMux I__7386 (
            .O(N__36640),
            .I(N__36634));
    LocalMux I__7385 (
            .O(N__36637),
            .I(N__36631));
    LocalMux I__7384 (
            .O(N__36634),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv12 I__7383 (
            .O(N__36631),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__7382 (
            .O(N__36626),
            .I(N__36623));
    InMux I__7381 (
            .O(N__36623),
            .I(N__36620));
    LocalMux I__7380 (
            .O(N__36620),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__7379 (
            .O(N__36617),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__7378 (
            .O(N__36614),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__7377 (
            .O(N__36611),
            .I(N__36605));
    InMux I__7376 (
            .O(N__36610),
            .I(N__36605));
    LocalMux I__7375 (
            .O(N__36605),
            .I(N__36602));
    Odrv12 I__7374 (
            .O(N__36602),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ));
    InMux I__7373 (
            .O(N__36599),
            .I(N__36594));
    InMux I__7372 (
            .O(N__36598),
            .I(N__36589));
    InMux I__7371 (
            .O(N__36597),
            .I(N__36589));
    LocalMux I__7370 (
            .O(N__36594),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__7369 (
            .O(N__36589),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    CascadeMux I__7368 (
            .O(N__36584),
            .I(N__36581));
    InMux I__7367 (
            .O(N__36581),
            .I(N__36574));
    InMux I__7366 (
            .O(N__36580),
            .I(N__36574));
    InMux I__7365 (
            .O(N__36579),
            .I(N__36571));
    LocalMux I__7364 (
            .O(N__36574),
            .I(N__36568));
    LocalMux I__7363 (
            .O(N__36571),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__7362 (
            .O(N__36568),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    CascadeMux I__7361 (
            .O(N__36563),
            .I(N__36560));
    InMux I__7360 (
            .O(N__36560),
            .I(N__36554));
    InMux I__7359 (
            .O(N__36559),
            .I(N__36554));
    LocalMux I__7358 (
            .O(N__36554),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ));
    CascadeMux I__7357 (
            .O(N__36551),
            .I(N__36548));
    InMux I__7356 (
            .O(N__36548),
            .I(N__36545));
    LocalMux I__7355 (
            .O(N__36545),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__7354 (
            .O(N__36542),
            .I(N__36539));
    LocalMux I__7353 (
            .O(N__36539),
            .I(N__36535));
    InMux I__7352 (
            .O(N__36538),
            .I(N__36532));
    Span4Mux_v I__7351 (
            .O(N__36535),
            .I(N__36529));
    LocalMux I__7350 (
            .O(N__36532),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__7349 (
            .O(N__36529),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__7348 (
            .O(N__36524),
            .I(N__36521));
    InMux I__7347 (
            .O(N__36521),
            .I(N__36518));
    LocalMux I__7346 (
            .O(N__36518),
            .I(N__36515));
    Odrv4 I__7345 (
            .O(N__36515),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__7344 (
            .O(N__36512),
            .I(N__36507));
    InMux I__7343 (
            .O(N__36511),
            .I(N__36504));
    InMux I__7342 (
            .O(N__36510),
            .I(N__36499));
    InMux I__7341 (
            .O(N__36507),
            .I(N__36499));
    LocalMux I__7340 (
            .O(N__36504),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    LocalMux I__7339 (
            .O(N__36499),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__7338 (
            .O(N__36494),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__7337 (
            .O(N__36491),
            .I(N__36486));
    InMux I__7336 (
            .O(N__36490),
            .I(N__36483));
    InMux I__7335 (
            .O(N__36489),
            .I(N__36478));
    InMux I__7334 (
            .O(N__36486),
            .I(N__36478));
    LocalMux I__7333 (
            .O(N__36483),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    LocalMux I__7332 (
            .O(N__36478),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__7331 (
            .O(N__36473),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    CascadeMux I__7330 (
            .O(N__36470),
            .I(N__36465));
    InMux I__7329 (
            .O(N__36469),
            .I(N__36462));
    InMux I__7328 (
            .O(N__36468),
            .I(N__36457));
    InMux I__7327 (
            .O(N__36465),
            .I(N__36457));
    LocalMux I__7326 (
            .O(N__36462),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    LocalMux I__7325 (
            .O(N__36457),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__7324 (
            .O(N__36452),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__7323 (
            .O(N__36449),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__7322 (
            .O(N__36446),
            .I(bfn_14_22_0_));
    InMux I__7321 (
            .O(N__36443),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__7320 (
            .O(N__36440),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__7319 (
            .O(N__36437),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__7318 (
            .O(N__36434),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__7317 (
            .O(N__36431),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__7316 (
            .O(N__36428),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__7315 (
            .O(N__36425),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__7314 (
            .O(N__36422),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__7313 (
            .O(N__36419),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__7312 (
            .O(N__36416),
            .I(bfn_14_21_0_));
    InMux I__7311 (
            .O(N__36413),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__7310 (
            .O(N__36410),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__7309 (
            .O(N__36407),
            .I(N__36402));
    InMux I__7308 (
            .O(N__36406),
            .I(N__36397));
    InMux I__7307 (
            .O(N__36405),
            .I(N__36397));
    LocalMux I__7306 (
            .O(N__36402),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    LocalMux I__7305 (
            .O(N__36397),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__7304 (
            .O(N__36392),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__7303 (
            .O(N__36389),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__7302 (
            .O(N__36386),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__7301 (
            .O(N__36383),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__7300 (
            .O(N__36380),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__7299 (
            .O(N__36377),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__7298 (
            .O(N__36374),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__7297 (
            .O(N__36371),
            .I(bfn_14_20_0_));
    InMux I__7296 (
            .O(N__36368),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__7295 (
            .O(N__36365),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    IoInMux I__7294 (
            .O(N__36362),
            .I(N__36359));
    LocalMux I__7293 (
            .O(N__36359),
            .I(N__36356));
    IoSpan4Mux I__7292 (
            .O(N__36356),
            .I(N__36353));
    Span4Mux_s3_v I__7291 (
            .O(N__36353),
            .I(N__36350));
    Sp12to4 I__7290 (
            .O(N__36350),
            .I(N__36347));
    Span12Mux_v I__7289 (
            .O(N__36347),
            .I(N__36344));
    Odrv12 I__7288 (
            .O(N__36344),
            .I(\pll_inst.red_c_i ));
    CascadeMux I__7287 (
            .O(N__36341),
            .I(N__36338));
    InMux I__7286 (
            .O(N__36338),
            .I(N__36333));
    InMux I__7285 (
            .O(N__36337),
            .I(N__36330));
    InMux I__7284 (
            .O(N__36336),
            .I(N__36327));
    LocalMux I__7283 (
            .O(N__36333),
            .I(N__36324));
    LocalMux I__7282 (
            .O(N__36330),
            .I(N__36321));
    LocalMux I__7281 (
            .O(N__36327),
            .I(N__36314));
    Span12Mux_h I__7280 (
            .O(N__36324),
            .I(N__36314));
    Sp12to4 I__7279 (
            .O(N__36321),
            .I(N__36314));
    Span12Mux_v I__7278 (
            .O(N__36314),
            .I(N__36311));
    Odrv12 I__7277 (
            .O(N__36311),
            .I(il_max_comp1_D2));
    InMux I__7276 (
            .O(N__36308),
            .I(N__36305));
    LocalMux I__7275 (
            .O(N__36305),
            .I(N__36301));
    InMux I__7274 (
            .O(N__36304),
            .I(N__36297));
    Span4Mux_v I__7273 (
            .O(N__36301),
            .I(N__36294));
    InMux I__7272 (
            .O(N__36300),
            .I(N__36291));
    LocalMux I__7271 (
            .O(N__36297),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    Odrv4 I__7270 (
            .O(N__36294),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    LocalMux I__7269 (
            .O(N__36291),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    InMux I__7268 (
            .O(N__36284),
            .I(N__36281));
    LocalMux I__7267 (
            .O(N__36281),
            .I(N__36277));
    InMux I__7266 (
            .O(N__36280),
            .I(N__36273));
    Span4Mux_v I__7265 (
            .O(N__36277),
            .I(N__36270));
    InMux I__7264 (
            .O(N__36276),
            .I(N__36267));
    LocalMux I__7263 (
            .O(N__36273),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv4 I__7262 (
            .O(N__36270),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    LocalMux I__7261 (
            .O(N__36267),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    InMux I__7260 (
            .O(N__36260),
            .I(N__36256));
    InMux I__7259 (
            .O(N__36259),
            .I(N__36252));
    LocalMux I__7258 (
            .O(N__36256),
            .I(N__36249));
    InMux I__7257 (
            .O(N__36255),
            .I(N__36246));
    LocalMux I__7256 (
            .O(N__36252),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    Odrv4 I__7255 (
            .O(N__36249),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    LocalMux I__7254 (
            .O(N__36246),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    InMux I__7253 (
            .O(N__36239),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__7252 (
            .O(N__36236),
            .I(N__36233));
    LocalMux I__7251 (
            .O(N__36233),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__7250 (
            .O(N__36230),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__7249 (
            .O(N__36227),
            .I(N__36224));
    LocalMux I__7248 (
            .O(N__36224),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__7247 (
            .O(N__36221),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__7246 (
            .O(N__36218),
            .I(N__36215));
    LocalMux I__7245 (
            .O(N__36215),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__7244 (
            .O(N__36212),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__7243 (
            .O(N__36209),
            .I(N__36206));
    LocalMux I__7242 (
            .O(N__36206),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__7241 (
            .O(N__36203),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__7240 (
            .O(N__36200),
            .I(N__36197));
    LocalMux I__7239 (
            .O(N__36197),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__7238 (
            .O(N__36194),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__7237 (
            .O(N__36191),
            .I(N__36188));
    LocalMux I__7236 (
            .O(N__36188),
            .I(N__36185));
    Odrv4 I__7235 (
            .O(N__36185),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__7234 (
            .O(N__36182),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    CascadeMux I__7233 (
            .O(N__36179),
            .I(N__36176));
    InMux I__7232 (
            .O(N__36176),
            .I(N__36173));
    LocalMux I__7231 (
            .O(N__36173),
            .I(N__36170));
    Span4Mux_v I__7230 (
            .O(N__36170),
            .I(N__36167));
    Odrv4 I__7229 (
            .O(N__36167),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__7228 (
            .O(N__36164),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__7227 (
            .O(N__36161),
            .I(N__36158));
    LocalMux I__7226 (
            .O(N__36158),
            .I(N__36155));
    Odrv4 I__7225 (
            .O(N__36155),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__7224 (
            .O(N__36152),
            .I(N__36149));
    LocalMux I__7223 (
            .O(N__36149),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__7222 (
            .O(N__36146),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__7221 (
            .O(N__36143),
            .I(N__36140));
    LocalMux I__7220 (
            .O(N__36140),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__7219 (
            .O(N__36137),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__7218 (
            .O(N__36134),
            .I(N__36131));
    LocalMux I__7217 (
            .O(N__36131),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__7216 (
            .O(N__36128),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__7215 (
            .O(N__36125),
            .I(N__36122));
    LocalMux I__7214 (
            .O(N__36122),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__7213 (
            .O(N__36119),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__7212 (
            .O(N__36116),
            .I(N__36113));
    LocalMux I__7211 (
            .O(N__36113),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__7210 (
            .O(N__36110),
            .I(bfn_14_12_0_));
    InMux I__7209 (
            .O(N__36107),
            .I(N__36104));
    LocalMux I__7208 (
            .O(N__36104),
            .I(N__36101));
    Odrv4 I__7207 (
            .O(N__36101),
            .I(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ));
    InMux I__7206 (
            .O(N__36098),
            .I(N__36095));
    LocalMux I__7205 (
            .O(N__36095),
            .I(N__36092));
    Span4Mux_v I__7204 (
            .O(N__36092),
            .I(N__36089));
    Odrv4 I__7203 (
            .O(N__36089),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__7202 (
            .O(N__36086),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__7201 (
            .O(N__36083),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__7200 (
            .O(N__36080),
            .I(N__36077));
    LocalMux I__7199 (
            .O(N__36077),
            .I(N__36074));
    Span4Mux_h I__7198 (
            .O(N__36074),
            .I(N__36071));
    Odrv4 I__7197 (
            .O(N__36071),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    CascadeMux I__7196 (
            .O(N__36068),
            .I(N__36065));
    InMux I__7195 (
            .O(N__36065),
            .I(N__36062));
    LocalMux I__7194 (
            .O(N__36062),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    CascadeMux I__7193 (
            .O(N__36059),
            .I(N__36056));
    InMux I__7192 (
            .O(N__36056),
            .I(N__36053));
    LocalMux I__7191 (
            .O(N__36053),
            .I(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ));
    InMux I__7190 (
            .O(N__36050),
            .I(N__36047));
    LocalMux I__7189 (
            .O(N__36047),
            .I(N__36044));
    Span4Mux_v I__7188 (
            .O(N__36044),
            .I(N__36041));
    Odrv4 I__7187 (
            .O(N__36041),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__7186 (
            .O(N__36038),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__7185 (
            .O(N__36035),
            .I(N__36032));
    LocalMux I__7184 (
            .O(N__36032),
            .I(N__36029));
    Span4Mux_v I__7183 (
            .O(N__36029),
            .I(N__36026));
    Odrv4 I__7182 (
            .O(N__36026),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__7181 (
            .O(N__36023),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    CascadeMux I__7180 (
            .O(N__36020),
            .I(N__36017));
    InMux I__7179 (
            .O(N__36017),
            .I(N__36014));
    LocalMux I__7178 (
            .O(N__36014),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__7177 (
            .O(N__36011),
            .I(N__36008));
    LocalMux I__7176 (
            .O(N__36008),
            .I(N__36005));
    Span4Mux_v I__7175 (
            .O(N__36005),
            .I(N__36002));
    Odrv4 I__7174 (
            .O(N__36002),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__7173 (
            .O(N__35999),
            .I(bfn_14_8_0_));
    InMux I__7172 (
            .O(N__35996),
            .I(N__35993));
    LocalMux I__7171 (
            .O(N__35993),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__7170 (
            .O(N__35990),
            .I(N__35987));
    LocalMux I__7169 (
            .O(N__35987),
            .I(N__35984));
    Span4Mux_v I__7168 (
            .O(N__35984),
            .I(N__35981));
    Odrv4 I__7167 (
            .O(N__35981),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__7166 (
            .O(N__35978),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    CascadeMux I__7165 (
            .O(N__35975),
            .I(N__35972));
    InMux I__7164 (
            .O(N__35972),
            .I(N__35969));
    LocalMux I__7163 (
            .O(N__35969),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__7162 (
            .O(N__35966),
            .I(N__35963));
    LocalMux I__7161 (
            .O(N__35963),
            .I(N__35960));
    Odrv4 I__7160 (
            .O(N__35960),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__7159 (
            .O(N__35957),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__7158 (
            .O(N__35954),
            .I(N__35951));
    LocalMux I__7157 (
            .O(N__35951),
            .I(N__35948));
    Odrv4 I__7156 (
            .O(N__35948),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__7155 (
            .O(N__35945),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__7154 (
            .O(N__35942),
            .I(N__35939));
    LocalMux I__7153 (
            .O(N__35939),
            .I(N__35936));
    Odrv4 I__7152 (
            .O(N__35936),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__7151 (
            .O(N__35933),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__7150 (
            .O(N__35930),
            .I(N__35927));
    LocalMux I__7149 (
            .O(N__35927),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__7148 (
            .O(N__35924),
            .I(N__35921));
    LocalMux I__7147 (
            .O(N__35921),
            .I(N__35918));
    Odrv4 I__7146 (
            .O(N__35918),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__7145 (
            .O(N__35915),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__7144 (
            .O(N__35912),
            .I(N__35909));
    LocalMux I__7143 (
            .O(N__35909),
            .I(N__35906));
    Span4Mux_h I__7142 (
            .O(N__35906),
            .I(N__35903));
    Odrv4 I__7141 (
            .O(N__35903),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__7140 (
            .O(N__35900),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__7139 (
            .O(N__35897),
            .I(N__35894));
    LocalMux I__7138 (
            .O(N__35894),
            .I(N__35891));
    Odrv4 I__7137 (
            .O(N__35891),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__7136 (
            .O(N__35888),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__7135 (
            .O(N__35885),
            .I(N__35882));
    LocalMux I__7134 (
            .O(N__35882),
            .I(N__35877));
    InMux I__7133 (
            .O(N__35881),
            .I(N__35874));
    InMux I__7132 (
            .O(N__35880),
            .I(N__35868));
    Span12Mux_h I__7131 (
            .O(N__35877),
            .I(N__35865));
    LocalMux I__7130 (
            .O(N__35874),
            .I(N__35862));
    InMux I__7129 (
            .O(N__35873),
            .I(N__35859));
    InMux I__7128 (
            .O(N__35872),
            .I(N__35856));
    InMux I__7127 (
            .O(N__35871),
            .I(N__35853));
    LocalMux I__7126 (
            .O(N__35868),
            .I(N__35850));
    Odrv12 I__7125 (
            .O(N__35865),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__7124 (
            .O(N__35862),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__7123 (
            .O(N__35859),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__7122 (
            .O(N__35856),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__7121 (
            .O(N__35853),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__7120 (
            .O(N__35850),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__7119 (
            .O(N__35837),
            .I(N__35834));
    LocalMux I__7118 (
            .O(N__35834),
            .I(N__35831));
    Odrv12 I__7117 (
            .O(N__35831),
            .I(s2_phy_c));
    CascadeMux I__7116 (
            .O(N__35828),
            .I(N__35825));
    InMux I__7115 (
            .O(N__35825),
            .I(N__35821));
    InMux I__7114 (
            .O(N__35824),
            .I(N__35818));
    LocalMux I__7113 (
            .O(N__35821),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    LocalMux I__7112 (
            .O(N__35818),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__7111 (
            .O(N__35813),
            .I(N__35808));
    InMux I__7110 (
            .O(N__35812),
            .I(N__35805));
    InMux I__7109 (
            .O(N__35811),
            .I(N__35801));
    LocalMux I__7108 (
            .O(N__35808),
            .I(N__35796));
    LocalMux I__7107 (
            .O(N__35805),
            .I(N__35796));
    CascadeMux I__7106 (
            .O(N__35804),
            .I(N__35793));
    LocalMux I__7105 (
            .O(N__35801),
            .I(N__35788));
    Span4Mux_v I__7104 (
            .O(N__35796),
            .I(N__35788));
    InMux I__7103 (
            .O(N__35793),
            .I(N__35785));
    Span4Mux_v I__7102 (
            .O(N__35788),
            .I(N__35782));
    LocalMux I__7101 (
            .O(N__35785),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__7100 (
            .O(N__35782),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    ClkMux I__7099 (
            .O(N__35777),
            .I(N__35774));
    GlobalMux I__7098 (
            .O(N__35774),
            .I(N__35771));
    gio2CtrlBuf I__7097 (
            .O(N__35771),
            .I(delay_hc_input_c_g));
    InMux I__7096 (
            .O(N__35768),
            .I(N__35765));
    LocalMux I__7095 (
            .O(N__35765),
            .I(N__35760));
    InMux I__7094 (
            .O(N__35764),
            .I(N__35757));
    InMux I__7093 (
            .O(N__35763),
            .I(N__35754));
    Span12Mux_v I__7092 (
            .O(N__35760),
            .I(N__35749));
    LocalMux I__7091 (
            .O(N__35757),
            .I(N__35749));
    LocalMux I__7090 (
            .O(N__35754),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    Odrv12 I__7089 (
            .O(N__35749),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    CascadeMux I__7088 (
            .O(N__35744),
            .I(N__35740));
    InMux I__7087 (
            .O(N__35743),
            .I(N__35736));
    InMux I__7086 (
            .O(N__35740),
            .I(N__35731));
    InMux I__7085 (
            .O(N__35739),
            .I(N__35731));
    LocalMux I__7084 (
            .O(N__35736),
            .I(N__35728));
    LocalMux I__7083 (
            .O(N__35731),
            .I(N__35725));
    Span12Mux_h I__7082 (
            .O(N__35728),
            .I(N__35721));
    Span12Mux_h I__7081 (
            .O(N__35725),
            .I(N__35718));
    InMux I__7080 (
            .O(N__35724),
            .I(N__35715));
    Span12Mux_v I__7079 (
            .O(N__35721),
            .I(N__35712));
    Span12Mux_v I__7078 (
            .O(N__35718),
            .I(N__35709));
    LocalMux I__7077 (
            .O(N__35715),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__7076 (
            .O(N__35712),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__7075 (
            .O(N__35709),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__7074 (
            .O(N__35702),
            .I(N__35696));
    InMux I__7073 (
            .O(N__35701),
            .I(N__35689));
    InMux I__7072 (
            .O(N__35700),
            .I(N__35689));
    InMux I__7071 (
            .O(N__35699),
            .I(N__35689));
    LocalMux I__7070 (
            .O(N__35696),
            .I(N__35686));
    LocalMux I__7069 (
            .O(N__35689),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv12 I__7068 (
            .O(N__35686),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    CascadeMux I__7067 (
            .O(N__35681),
            .I(N__35676));
    InMux I__7066 (
            .O(N__35680),
            .I(N__35672));
    InMux I__7065 (
            .O(N__35679),
            .I(N__35669));
    InMux I__7064 (
            .O(N__35676),
            .I(N__35664));
    InMux I__7063 (
            .O(N__35675),
            .I(N__35664));
    LocalMux I__7062 (
            .O(N__35672),
            .I(N__35661));
    LocalMux I__7061 (
            .O(N__35669),
            .I(N__35658));
    LocalMux I__7060 (
            .O(N__35664),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv12 I__7059 (
            .O(N__35661),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv4 I__7058 (
            .O(N__35658),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    InMux I__7057 (
            .O(N__35651),
            .I(N__35647));
    InMux I__7056 (
            .O(N__35650),
            .I(N__35642));
    LocalMux I__7055 (
            .O(N__35647),
            .I(N__35639));
    InMux I__7054 (
            .O(N__35646),
            .I(N__35636));
    InMux I__7053 (
            .O(N__35645),
            .I(N__35633));
    LocalMux I__7052 (
            .O(N__35642),
            .I(N__35628));
    Span12Mux_v I__7051 (
            .O(N__35639),
            .I(N__35628));
    LocalMux I__7050 (
            .O(N__35636),
            .I(N__35625));
    LocalMux I__7049 (
            .O(N__35633),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__7048 (
            .O(N__35628),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__7047 (
            .O(N__35625),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    IoInMux I__7046 (
            .O(N__35618),
            .I(N__35615));
    LocalMux I__7045 (
            .O(N__35615),
            .I(N__35612));
    Span4Mux_s1_v I__7044 (
            .O(N__35612),
            .I(N__35609));
    Span4Mux_v I__7043 (
            .O(N__35609),
            .I(N__35604));
    InMux I__7042 (
            .O(N__35608),
            .I(N__35599));
    InMux I__7041 (
            .O(N__35607),
            .I(N__35599));
    Odrv4 I__7040 (
            .O(N__35604),
            .I(s1_phy_c));
    LocalMux I__7039 (
            .O(N__35599),
            .I(s1_phy_c));
    InMux I__7038 (
            .O(N__35594),
            .I(N__35591));
    LocalMux I__7037 (
            .O(N__35591),
            .I(N__35588));
    Odrv12 I__7036 (
            .O(N__35588),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    CascadeMux I__7035 (
            .O(N__35585),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    IoInMux I__7034 (
            .O(N__35582),
            .I(N__35579));
    LocalMux I__7033 (
            .O(N__35579),
            .I(N__35576));
    Odrv12 I__7032 (
            .O(N__35576),
            .I(\current_shift_inst.timer_s1.N_167_i ));
    InMux I__7031 (
            .O(N__35573),
            .I(N__35570));
    LocalMux I__7030 (
            .O(N__35570),
            .I(N__35565));
    InMux I__7029 (
            .O(N__35569),
            .I(N__35562));
    InMux I__7028 (
            .O(N__35568),
            .I(N__35559));
    Span4Mux_v I__7027 (
            .O(N__35565),
            .I(N__35554));
    LocalMux I__7026 (
            .O(N__35562),
            .I(N__35554));
    LocalMux I__7025 (
            .O(N__35559),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    Odrv4 I__7024 (
            .O(N__35554),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    InMux I__7023 (
            .O(N__35549),
            .I(N__35543));
    InMux I__7022 (
            .O(N__35548),
            .I(N__35543));
    LocalMux I__7021 (
            .O(N__35543),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    InMux I__7020 (
            .O(N__35540),
            .I(N__35534));
    InMux I__7019 (
            .O(N__35539),
            .I(N__35534));
    LocalMux I__7018 (
            .O(N__35534),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    InMux I__7017 (
            .O(N__35531),
            .I(N__35525));
    InMux I__7016 (
            .O(N__35530),
            .I(N__35525));
    LocalMux I__7015 (
            .O(N__35525),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ));
    CascadeMux I__7014 (
            .O(N__35522),
            .I(N__35519));
    InMux I__7013 (
            .O(N__35519),
            .I(N__35513));
    InMux I__7012 (
            .O(N__35518),
            .I(N__35513));
    LocalMux I__7011 (
            .O(N__35513),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ));
    IoInMux I__7010 (
            .O(N__35510),
            .I(N__35507));
    LocalMux I__7009 (
            .O(N__35507),
            .I(N__35504));
    Span4Mux_s2_v I__7008 (
            .O(N__35504),
            .I(N__35501));
    Span4Mux_h I__7007 (
            .O(N__35501),
            .I(N__35498));
    Span4Mux_v I__7006 (
            .O(N__35498),
            .I(N__35495));
    Span4Mux_v I__7005 (
            .O(N__35495),
            .I(N__35491));
    InMux I__7004 (
            .O(N__35494),
            .I(N__35488));
    Odrv4 I__7003 (
            .O(N__35491),
            .I(T12_c));
    LocalMux I__7002 (
            .O(N__35488),
            .I(T12_c));
    CascadeMux I__7001 (
            .O(N__35483),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_ ));
    InMux I__7000 (
            .O(N__35480),
            .I(N__35477));
    LocalMux I__6999 (
            .O(N__35477),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ));
    CascadeMux I__6998 (
            .O(N__35474),
            .I(N__35468));
    CascadeMux I__6997 (
            .O(N__35473),
            .I(N__35465));
    InMux I__6996 (
            .O(N__35472),
            .I(N__35462));
    InMux I__6995 (
            .O(N__35471),
            .I(N__35458));
    InMux I__6994 (
            .O(N__35468),
            .I(N__35453));
    InMux I__6993 (
            .O(N__35465),
            .I(N__35453));
    LocalMux I__6992 (
            .O(N__35462),
            .I(N__35450));
    InMux I__6991 (
            .O(N__35461),
            .I(N__35447));
    LocalMux I__6990 (
            .O(N__35458),
            .I(N__35444));
    LocalMux I__6989 (
            .O(N__35453),
            .I(N__35441));
    Span4Mux_h I__6988 (
            .O(N__35450),
            .I(N__35438));
    LocalMux I__6987 (
            .O(N__35447),
            .I(N__35435));
    Span4Mux_h I__6986 (
            .O(N__35444),
            .I(N__35432));
    Span4Mux_v I__6985 (
            .O(N__35441),
            .I(N__35427));
    Span4Mux_v I__6984 (
            .O(N__35438),
            .I(N__35427));
    Odrv4 I__6983 (
            .O(N__35435),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__6982 (
            .O(N__35432),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__6981 (
            .O(N__35427),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__6980 (
            .O(N__35420),
            .I(N__35417));
    LocalMux I__6979 (
            .O(N__35417),
            .I(N__35414));
    Span4Mux_h I__6978 (
            .O(N__35414),
            .I(N__35411));
    Span4Mux_h I__6977 (
            .O(N__35411),
            .I(N__35408));
    Odrv4 I__6976 (
            .O(N__35408),
            .I(\current_shift_inst.PI_CTRL.integrator_i_19 ));
    CascadeMux I__6975 (
            .O(N__35405),
            .I(N__35392));
    CascadeMux I__6974 (
            .O(N__35404),
            .I(N__35388));
    CascadeMux I__6973 (
            .O(N__35403),
            .I(N__35385));
    InMux I__6972 (
            .O(N__35402),
            .I(N__35377));
    CascadeMux I__6971 (
            .O(N__35401),
            .I(N__35372));
    CascadeMux I__6970 (
            .O(N__35400),
            .I(N__35369));
    CascadeMux I__6969 (
            .O(N__35399),
            .I(N__35365));
    CascadeMux I__6968 (
            .O(N__35398),
            .I(N__35362));
    CascadeMux I__6967 (
            .O(N__35397),
            .I(N__35359));
    CascadeMux I__6966 (
            .O(N__35396),
            .I(N__35355));
    CascadeMux I__6965 (
            .O(N__35395),
            .I(N__35351));
    InMux I__6964 (
            .O(N__35392),
            .I(N__35348));
    InMux I__6963 (
            .O(N__35391),
            .I(N__35343));
    InMux I__6962 (
            .O(N__35388),
            .I(N__35343));
    InMux I__6961 (
            .O(N__35385),
            .I(N__35340));
    CascadeMux I__6960 (
            .O(N__35384),
            .I(N__35327));
    CascadeMux I__6959 (
            .O(N__35383),
            .I(N__35324));
    CascadeMux I__6958 (
            .O(N__35382),
            .I(N__35321));
    CascadeMux I__6957 (
            .O(N__35381),
            .I(N__35317));
    CascadeMux I__6956 (
            .O(N__35380),
            .I(N__35314));
    LocalMux I__6955 (
            .O(N__35377),
            .I(N__35311));
    InMux I__6954 (
            .O(N__35376),
            .I(N__35302));
    InMux I__6953 (
            .O(N__35375),
            .I(N__35302));
    InMux I__6952 (
            .O(N__35372),
            .I(N__35302));
    InMux I__6951 (
            .O(N__35369),
            .I(N__35302));
    InMux I__6950 (
            .O(N__35368),
            .I(N__35293));
    InMux I__6949 (
            .O(N__35365),
            .I(N__35293));
    InMux I__6948 (
            .O(N__35362),
            .I(N__35293));
    InMux I__6947 (
            .O(N__35359),
            .I(N__35293));
    InMux I__6946 (
            .O(N__35358),
            .I(N__35289));
    InMux I__6945 (
            .O(N__35355),
            .I(N__35282));
    InMux I__6944 (
            .O(N__35354),
            .I(N__35282));
    InMux I__6943 (
            .O(N__35351),
            .I(N__35282));
    LocalMux I__6942 (
            .O(N__35348),
            .I(N__35279));
    LocalMux I__6941 (
            .O(N__35343),
            .I(N__35274));
    LocalMux I__6940 (
            .O(N__35340),
            .I(N__35274));
    InMux I__6939 (
            .O(N__35339),
            .I(N__35261));
    InMux I__6938 (
            .O(N__35338),
            .I(N__35261));
    InMux I__6937 (
            .O(N__35337),
            .I(N__35261));
    InMux I__6936 (
            .O(N__35336),
            .I(N__35261));
    InMux I__6935 (
            .O(N__35335),
            .I(N__35261));
    InMux I__6934 (
            .O(N__35334),
            .I(N__35261));
    InMux I__6933 (
            .O(N__35333),
            .I(N__35254));
    InMux I__6932 (
            .O(N__35332),
            .I(N__35254));
    InMux I__6931 (
            .O(N__35331),
            .I(N__35254));
    InMux I__6930 (
            .O(N__35330),
            .I(N__35240));
    InMux I__6929 (
            .O(N__35327),
            .I(N__35240));
    InMux I__6928 (
            .O(N__35324),
            .I(N__35240));
    InMux I__6927 (
            .O(N__35321),
            .I(N__35240));
    InMux I__6926 (
            .O(N__35320),
            .I(N__35240));
    InMux I__6925 (
            .O(N__35317),
            .I(N__35240));
    InMux I__6924 (
            .O(N__35314),
            .I(N__35228));
    Span4Mux_v I__6923 (
            .O(N__35311),
            .I(N__35221));
    LocalMux I__6922 (
            .O(N__35302),
            .I(N__35221));
    LocalMux I__6921 (
            .O(N__35293),
            .I(N__35221));
    InMux I__6920 (
            .O(N__35292),
            .I(N__35218));
    LocalMux I__6919 (
            .O(N__35289),
            .I(N__35204));
    LocalMux I__6918 (
            .O(N__35282),
            .I(N__35204));
    Span4Mux_h I__6917 (
            .O(N__35279),
            .I(N__35204));
    Span4Mux_v I__6916 (
            .O(N__35274),
            .I(N__35204));
    LocalMux I__6915 (
            .O(N__35261),
            .I(N__35204));
    LocalMux I__6914 (
            .O(N__35254),
            .I(N__35204));
    InMux I__6913 (
            .O(N__35253),
            .I(N__35201));
    LocalMux I__6912 (
            .O(N__35240),
            .I(N__35198));
    InMux I__6911 (
            .O(N__35239),
            .I(N__35195));
    InMux I__6910 (
            .O(N__35238),
            .I(N__35178));
    InMux I__6909 (
            .O(N__35237),
            .I(N__35178));
    InMux I__6908 (
            .O(N__35236),
            .I(N__35178));
    InMux I__6907 (
            .O(N__35235),
            .I(N__35178));
    InMux I__6906 (
            .O(N__35234),
            .I(N__35178));
    InMux I__6905 (
            .O(N__35233),
            .I(N__35178));
    InMux I__6904 (
            .O(N__35232),
            .I(N__35178));
    InMux I__6903 (
            .O(N__35231),
            .I(N__35178));
    LocalMux I__6902 (
            .O(N__35228),
            .I(N__35171));
    Span4Mux_v I__6901 (
            .O(N__35221),
            .I(N__35166));
    LocalMux I__6900 (
            .O(N__35218),
            .I(N__35166));
    InMux I__6899 (
            .O(N__35217),
            .I(N__35163));
    Span4Mux_v I__6898 (
            .O(N__35204),
            .I(N__35160));
    LocalMux I__6897 (
            .O(N__35201),
            .I(N__35151));
    Span4Mux_h I__6896 (
            .O(N__35198),
            .I(N__35151));
    LocalMux I__6895 (
            .O(N__35195),
            .I(N__35151));
    LocalMux I__6894 (
            .O(N__35178),
            .I(N__35151));
    InMux I__6893 (
            .O(N__35177),
            .I(N__35142));
    InMux I__6892 (
            .O(N__35176),
            .I(N__35142));
    InMux I__6891 (
            .O(N__35175),
            .I(N__35142));
    InMux I__6890 (
            .O(N__35174),
            .I(N__35142));
    Odrv12 I__6889 (
            .O(N__35171),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__6888 (
            .O(N__35166),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    LocalMux I__6887 (
            .O(N__35163),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__6886 (
            .O(N__35160),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__6885 (
            .O(N__35151),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    LocalMux I__6884 (
            .O(N__35142),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__6883 (
            .O(N__35129),
            .I(N__35125));
    InMux I__6882 (
            .O(N__35128),
            .I(N__35122));
    LocalMux I__6881 (
            .O(N__35125),
            .I(N__35116));
    LocalMux I__6880 (
            .O(N__35122),
            .I(N__35116));
    InMux I__6879 (
            .O(N__35121),
            .I(N__35113));
    Span4Mux_h I__6878 (
            .O(N__35116),
            .I(N__35110));
    LocalMux I__6877 (
            .O(N__35113),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv4 I__6876 (
            .O(N__35110),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    InMux I__6875 (
            .O(N__35105),
            .I(N__35102));
    LocalMux I__6874 (
            .O(N__35102),
            .I(\phase_controller_inst1.N_55 ));
    InMux I__6873 (
            .O(N__35099),
            .I(N__35093));
    InMux I__6872 (
            .O(N__35098),
            .I(N__35093));
    LocalMux I__6871 (
            .O(N__35093),
            .I(N__35089));
    InMux I__6870 (
            .O(N__35092),
            .I(N__35085));
    Span4Mux_h I__6869 (
            .O(N__35089),
            .I(N__35082));
    InMux I__6868 (
            .O(N__35088),
            .I(N__35079));
    LocalMux I__6867 (
            .O(N__35085),
            .I(N__35076));
    Span4Mux_v I__6866 (
            .O(N__35082),
            .I(N__35073));
    LocalMux I__6865 (
            .O(N__35079),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__6864 (
            .O(N__35076),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__6863 (
            .O(N__35073),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__6862 (
            .O(N__35066),
            .I(N__35062));
    InMux I__6861 (
            .O(N__35065),
            .I(N__35059));
    LocalMux I__6860 (
            .O(N__35062),
            .I(N__35053));
    LocalMux I__6859 (
            .O(N__35059),
            .I(N__35053));
    InMux I__6858 (
            .O(N__35058),
            .I(N__35050));
    Span4Mux_s3_v I__6857 (
            .O(N__35053),
            .I(N__35047));
    LocalMux I__6856 (
            .O(N__35050),
            .I(N__35044));
    Span4Mux_h I__6855 (
            .O(N__35047),
            .I(N__35041));
    Span4Mux_v I__6854 (
            .O(N__35044),
            .I(N__35038));
    Sp12to4 I__6853 (
            .O(N__35041),
            .I(N__35034));
    Span4Mux_h I__6852 (
            .O(N__35038),
            .I(N__35031));
    InMux I__6851 (
            .O(N__35037),
            .I(N__35028));
    Span12Mux_v I__6850 (
            .O(N__35034),
            .I(N__35025));
    Sp12to4 I__6849 (
            .O(N__35031),
            .I(N__35022));
    LocalMux I__6848 (
            .O(N__35028),
            .I(N__35019));
    Span12Mux_v I__6847 (
            .O(N__35025),
            .I(N__35016));
    Span12Mux_s7_h I__6846 (
            .O(N__35022),
            .I(N__35011));
    Span12Mux_h I__6845 (
            .O(N__35019),
            .I(N__35011));
    Span12Mux_h I__6844 (
            .O(N__35016),
            .I(N__35006));
    Span12Mux_v I__6843 (
            .O(N__35011),
            .I(N__35006));
    Odrv12 I__6842 (
            .O(N__35006),
            .I(start_stop_c));
    InMux I__6841 (
            .O(N__35003),
            .I(N__34999));
    InMux I__6840 (
            .O(N__35002),
            .I(N__34996));
    LocalMux I__6839 (
            .O(N__34999),
            .I(N__34993));
    LocalMux I__6838 (
            .O(N__34996),
            .I(N__34990));
    Span12Mux_s9_v I__6837 (
            .O(N__34993),
            .I(N__34987));
    Odrv4 I__6836 (
            .O(N__34990),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv12 I__6835 (
            .O(N__34987),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    CascadeMux I__6834 (
            .O(N__34982),
            .I(N__34979));
    InMux I__6833 (
            .O(N__34979),
            .I(N__34976));
    LocalMux I__6832 (
            .O(N__34976),
            .I(N__34972));
    InMux I__6831 (
            .O(N__34975),
            .I(N__34969));
    Span4Mux_v I__6830 (
            .O(N__34972),
            .I(N__34966));
    LocalMux I__6829 (
            .O(N__34969),
            .I(N__34963));
    Span4Mux_v I__6828 (
            .O(N__34966),
            .I(N__34955));
    Span4Mux_v I__6827 (
            .O(N__34963),
            .I(N__34955));
    InMux I__6826 (
            .O(N__34962),
            .I(N__34948));
    InMux I__6825 (
            .O(N__34961),
            .I(N__34948));
    InMux I__6824 (
            .O(N__34960),
            .I(N__34948));
    Odrv4 I__6823 (
            .O(N__34955),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__6822 (
            .O(N__34948),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__6821 (
            .O(N__34943),
            .I(N__34938));
    InMux I__6820 (
            .O(N__34942),
            .I(N__34935));
    CascadeMux I__6819 (
            .O(N__34941),
            .I(N__34932));
    LocalMux I__6818 (
            .O(N__34938),
            .I(N__34929));
    LocalMux I__6817 (
            .O(N__34935),
            .I(N__34926));
    InMux I__6816 (
            .O(N__34932),
            .I(N__34922));
    Span4Mux_v I__6815 (
            .O(N__34929),
            .I(N__34919));
    Span12Mux_v I__6814 (
            .O(N__34926),
            .I(N__34916));
    InMux I__6813 (
            .O(N__34925),
            .I(N__34913));
    LocalMux I__6812 (
            .O(N__34922),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv4 I__6811 (
            .O(N__34919),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv12 I__6810 (
            .O(N__34916),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__6809 (
            .O(N__34913),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__6808 (
            .O(N__34904),
            .I(N__34899));
    InMux I__6807 (
            .O(N__34903),
            .I(N__34894));
    InMux I__6806 (
            .O(N__34902),
            .I(N__34894));
    LocalMux I__6805 (
            .O(N__34899),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__6804 (
            .O(N__34894),
            .I(\phase_controller_inst1.tr_time_passed ));
    CascadeMux I__6803 (
            .O(N__34889),
            .I(N__34885));
    CascadeMux I__6802 (
            .O(N__34888),
            .I(N__34881));
    InMux I__6801 (
            .O(N__34885),
            .I(N__34878));
    InMux I__6800 (
            .O(N__34884),
            .I(N__34875));
    InMux I__6799 (
            .O(N__34881),
            .I(N__34872));
    LocalMux I__6798 (
            .O(N__34878),
            .I(N__34869));
    LocalMux I__6797 (
            .O(N__34875),
            .I(N__34864));
    LocalMux I__6796 (
            .O(N__34872),
            .I(N__34864));
    Span12Mux_h I__6795 (
            .O(N__34869),
            .I(N__34861));
    Span12Mux_v I__6794 (
            .O(N__34864),
            .I(N__34858));
    Span12Mux_v I__6793 (
            .O(N__34861),
            .I(N__34855));
    Odrv12 I__6792 (
            .O(N__34858),
            .I(il_min_comp1_D2));
    Odrv12 I__6791 (
            .O(N__34855),
            .I(il_min_comp1_D2));
    CascadeMux I__6790 (
            .O(N__34850),
            .I(N__34847));
    InMux I__6789 (
            .O(N__34847),
            .I(N__34844));
    LocalMux I__6788 (
            .O(N__34844),
            .I(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ));
    InMux I__6787 (
            .O(N__34841),
            .I(N__34838));
    LocalMux I__6786 (
            .O(N__34838),
            .I(N__34833));
    InMux I__6785 (
            .O(N__34837),
            .I(N__34830));
    InMux I__6784 (
            .O(N__34836),
            .I(N__34827));
    Span4Mux_v I__6783 (
            .O(N__34833),
            .I(N__34824));
    LocalMux I__6782 (
            .O(N__34830),
            .I(N__34821));
    LocalMux I__6781 (
            .O(N__34827),
            .I(N__34811));
    Span4Mux_h I__6780 (
            .O(N__34824),
            .I(N__34811));
    Span4Mux_h I__6779 (
            .O(N__34821),
            .I(N__34811));
    InMux I__6778 (
            .O(N__34820),
            .I(N__34806));
    InMux I__6777 (
            .O(N__34819),
            .I(N__34806));
    InMux I__6776 (
            .O(N__34818),
            .I(N__34803));
    Odrv4 I__6775 (
            .O(N__34811),
            .I(phase_controller_inst1_state_4));
    LocalMux I__6774 (
            .O(N__34806),
            .I(phase_controller_inst1_state_4));
    LocalMux I__6773 (
            .O(N__34803),
            .I(phase_controller_inst1_state_4));
    InMux I__6772 (
            .O(N__34796),
            .I(N__34793));
    LocalMux I__6771 (
            .O(N__34793),
            .I(N__34789));
    InMux I__6770 (
            .O(N__34792),
            .I(N__34786));
    Odrv4 I__6769 (
            .O(N__34789),
            .I(\phase_controller_inst1.N_54 ));
    LocalMux I__6768 (
            .O(N__34786),
            .I(\phase_controller_inst1.N_54 ));
    CascadeMux I__6767 (
            .O(N__34781),
            .I(N__34778));
    InMux I__6766 (
            .O(N__34778),
            .I(N__34775));
    LocalMux I__6765 (
            .O(N__34775),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__6764 (
            .O(N__34772),
            .I(N__34769));
    LocalMux I__6763 (
            .O(N__34769),
            .I(N__34764));
    InMux I__6762 (
            .O(N__34768),
            .I(N__34761));
    InMux I__6761 (
            .O(N__34767),
            .I(N__34758));
    Span4Mux_v I__6760 (
            .O(N__34764),
            .I(N__34755));
    LocalMux I__6759 (
            .O(N__34761),
            .I(N__34752));
    LocalMux I__6758 (
            .O(N__34758),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    Odrv4 I__6757 (
            .O(N__34755),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    Odrv12 I__6756 (
            .O(N__34752),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    InMux I__6755 (
            .O(N__34745),
            .I(N__34740));
    InMux I__6754 (
            .O(N__34744),
            .I(N__34737));
    InMux I__6753 (
            .O(N__34743),
            .I(N__34734));
    LocalMux I__6752 (
            .O(N__34740),
            .I(N__34731));
    LocalMux I__6751 (
            .O(N__34737),
            .I(N__34728));
    LocalMux I__6750 (
            .O(N__34734),
            .I(N__34725));
    Span4Mux_v I__6749 (
            .O(N__34731),
            .I(N__34721));
    Span4Mux_v I__6748 (
            .O(N__34728),
            .I(N__34716));
    Span4Mux_v I__6747 (
            .O(N__34725),
            .I(N__34716));
    InMux I__6746 (
            .O(N__34724),
            .I(N__34713));
    Odrv4 I__6745 (
            .O(N__34721),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv4 I__6744 (
            .O(N__34716),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__6743 (
            .O(N__34713),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    CascadeMux I__6742 (
            .O(N__34706),
            .I(N__34690));
    CascadeMux I__6741 (
            .O(N__34705),
            .I(N__34669));
    InMux I__6740 (
            .O(N__34704),
            .I(N__34651));
    InMux I__6739 (
            .O(N__34703),
            .I(N__34651));
    InMux I__6738 (
            .O(N__34702),
            .I(N__34651));
    InMux I__6737 (
            .O(N__34701),
            .I(N__34651));
    InMux I__6736 (
            .O(N__34700),
            .I(N__34651));
    InMux I__6735 (
            .O(N__34699),
            .I(N__34642));
    InMux I__6734 (
            .O(N__34698),
            .I(N__34642));
    InMux I__6733 (
            .O(N__34697),
            .I(N__34642));
    InMux I__6732 (
            .O(N__34696),
            .I(N__34642));
    InMux I__6731 (
            .O(N__34695),
            .I(N__34629));
    InMux I__6730 (
            .O(N__34694),
            .I(N__34629));
    InMux I__6729 (
            .O(N__34693),
            .I(N__34629));
    InMux I__6728 (
            .O(N__34690),
            .I(N__34629));
    InMux I__6727 (
            .O(N__34689),
            .I(N__34629));
    InMux I__6726 (
            .O(N__34688),
            .I(N__34629));
    InMux I__6725 (
            .O(N__34687),
            .I(N__34626));
    InMux I__6724 (
            .O(N__34686),
            .I(N__34617));
    InMux I__6723 (
            .O(N__34685),
            .I(N__34617));
    CascadeMux I__6722 (
            .O(N__34684),
            .I(N__34599));
    InMux I__6721 (
            .O(N__34683),
            .I(N__34579));
    InMux I__6720 (
            .O(N__34682),
            .I(N__34579));
    InMux I__6719 (
            .O(N__34681),
            .I(N__34579));
    InMux I__6718 (
            .O(N__34680),
            .I(N__34562));
    InMux I__6717 (
            .O(N__34679),
            .I(N__34562));
    InMux I__6716 (
            .O(N__34678),
            .I(N__34562));
    InMux I__6715 (
            .O(N__34677),
            .I(N__34562));
    InMux I__6714 (
            .O(N__34676),
            .I(N__34562));
    InMux I__6713 (
            .O(N__34675),
            .I(N__34562));
    InMux I__6712 (
            .O(N__34674),
            .I(N__34551));
    InMux I__6711 (
            .O(N__34673),
            .I(N__34551));
    InMux I__6710 (
            .O(N__34672),
            .I(N__34551));
    InMux I__6709 (
            .O(N__34669),
            .I(N__34551));
    InMux I__6708 (
            .O(N__34668),
            .I(N__34551));
    InMux I__6707 (
            .O(N__34667),
            .I(N__34538));
    InMux I__6706 (
            .O(N__34666),
            .I(N__34538));
    InMux I__6705 (
            .O(N__34665),
            .I(N__34538));
    InMux I__6704 (
            .O(N__34664),
            .I(N__34538));
    InMux I__6703 (
            .O(N__34663),
            .I(N__34538));
    InMux I__6702 (
            .O(N__34662),
            .I(N__34538));
    LocalMux I__6701 (
            .O(N__34651),
            .I(N__34533));
    LocalMux I__6700 (
            .O(N__34642),
            .I(N__34533));
    LocalMux I__6699 (
            .O(N__34629),
            .I(N__34529));
    LocalMux I__6698 (
            .O(N__34626),
            .I(N__34526));
    InMux I__6697 (
            .O(N__34625),
            .I(N__34521));
    InMux I__6696 (
            .O(N__34624),
            .I(N__34521));
    InMux I__6695 (
            .O(N__34623),
            .I(N__34516));
    InMux I__6694 (
            .O(N__34622),
            .I(N__34516));
    LocalMux I__6693 (
            .O(N__34617),
            .I(N__34508));
    InMux I__6692 (
            .O(N__34616),
            .I(N__34501));
    InMux I__6691 (
            .O(N__34615),
            .I(N__34501));
    InMux I__6690 (
            .O(N__34614),
            .I(N__34501));
    InMux I__6689 (
            .O(N__34613),
            .I(N__34496));
    InMux I__6688 (
            .O(N__34612),
            .I(N__34496));
    InMux I__6687 (
            .O(N__34611),
            .I(N__34491));
    InMux I__6686 (
            .O(N__34610),
            .I(N__34491));
    InMux I__6685 (
            .O(N__34609),
            .I(N__34488));
    InMux I__6684 (
            .O(N__34608),
            .I(N__34485));
    CascadeMux I__6683 (
            .O(N__34607),
            .I(N__34477));
    InMux I__6682 (
            .O(N__34606),
            .I(N__34473));
    InMux I__6681 (
            .O(N__34605),
            .I(N__34457));
    InMux I__6680 (
            .O(N__34604),
            .I(N__34457));
    InMux I__6679 (
            .O(N__34603),
            .I(N__34457));
    InMux I__6678 (
            .O(N__34602),
            .I(N__34457));
    InMux I__6677 (
            .O(N__34599),
            .I(N__34457));
    InMux I__6676 (
            .O(N__34598),
            .I(N__34454));
    InMux I__6675 (
            .O(N__34597),
            .I(N__34441));
    InMux I__6674 (
            .O(N__34596),
            .I(N__34441));
    InMux I__6673 (
            .O(N__34595),
            .I(N__34441));
    InMux I__6672 (
            .O(N__34594),
            .I(N__34441));
    InMux I__6671 (
            .O(N__34593),
            .I(N__34441));
    InMux I__6670 (
            .O(N__34592),
            .I(N__34441));
    InMux I__6669 (
            .O(N__34591),
            .I(N__34430));
    InMux I__6668 (
            .O(N__34590),
            .I(N__34430));
    InMux I__6667 (
            .O(N__34589),
            .I(N__34430));
    InMux I__6666 (
            .O(N__34588),
            .I(N__34430));
    InMux I__6665 (
            .O(N__34587),
            .I(N__34430));
    InMux I__6664 (
            .O(N__34586),
            .I(N__34427));
    LocalMux I__6663 (
            .O(N__34579),
            .I(N__34424));
    InMux I__6662 (
            .O(N__34578),
            .I(N__34415));
    InMux I__6661 (
            .O(N__34577),
            .I(N__34415));
    InMux I__6660 (
            .O(N__34576),
            .I(N__34415));
    InMux I__6659 (
            .O(N__34575),
            .I(N__34415));
    LocalMux I__6658 (
            .O(N__34562),
            .I(N__34406));
    LocalMux I__6657 (
            .O(N__34551),
            .I(N__34406));
    LocalMux I__6656 (
            .O(N__34538),
            .I(N__34406));
    Span4Mux_v I__6655 (
            .O(N__34533),
            .I(N__34406));
    InMux I__6654 (
            .O(N__34532),
            .I(N__34403));
    Span4Mux_h I__6653 (
            .O(N__34529),
            .I(N__34396));
    Span4Mux_v I__6652 (
            .O(N__34526),
            .I(N__34396));
    LocalMux I__6651 (
            .O(N__34521),
            .I(N__34396));
    LocalMux I__6650 (
            .O(N__34516),
            .I(N__34393));
    InMux I__6649 (
            .O(N__34515),
            .I(N__34382));
    InMux I__6648 (
            .O(N__34514),
            .I(N__34382));
    InMux I__6647 (
            .O(N__34513),
            .I(N__34382));
    InMux I__6646 (
            .O(N__34512),
            .I(N__34382));
    InMux I__6645 (
            .O(N__34511),
            .I(N__34382));
    Span4Mux_v I__6644 (
            .O(N__34508),
            .I(N__34377));
    LocalMux I__6643 (
            .O(N__34501),
            .I(N__34377));
    LocalMux I__6642 (
            .O(N__34496),
            .I(N__34372));
    LocalMux I__6641 (
            .O(N__34491),
            .I(N__34372));
    LocalMux I__6640 (
            .O(N__34488),
            .I(N__34369));
    LocalMux I__6639 (
            .O(N__34485),
            .I(N__34366));
    InMux I__6638 (
            .O(N__34484),
            .I(N__34359));
    InMux I__6637 (
            .O(N__34483),
            .I(N__34359));
    InMux I__6636 (
            .O(N__34482),
            .I(N__34359));
    InMux I__6635 (
            .O(N__34481),
            .I(N__34354));
    InMux I__6634 (
            .O(N__34480),
            .I(N__34354));
    InMux I__6633 (
            .O(N__34477),
            .I(N__34349));
    InMux I__6632 (
            .O(N__34476),
            .I(N__34349));
    LocalMux I__6631 (
            .O(N__34473),
            .I(N__34346));
    InMux I__6630 (
            .O(N__34472),
            .I(N__34335));
    InMux I__6629 (
            .O(N__34471),
            .I(N__34335));
    InMux I__6628 (
            .O(N__34470),
            .I(N__34335));
    InMux I__6627 (
            .O(N__34469),
            .I(N__34335));
    InMux I__6626 (
            .O(N__34468),
            .I(N__34335));
    LocalMux I__6625 (
            .O(N__34457),
            .I(N__34326));
    LocalMux I__6624 (
            .O(N__34454),
            .I(N__34326));
    LocalMux I__6623 (
            .O(N__34441),
            .I(N__34326));
    LocalMux I__6622 (
            .O(N__34430),
            .I(N__34326));
    LocalMux I__6621 (
            .O(N__34427),
            .I(N__34317));
    Span4Mux_v I__6620 (
            .O(N__34424),
            .I(N__34317));
    LocalMux I__6619 (
            .O(N__34415),
            .I(N__34317));
    Span4Mux_v I__6618 (
            .O(N__34406),
            .I(N__34317));
    LocalMux I__6617 (
            .O(N__34403),
            .I(N__34312));
    Span4Mux_h I__6616 (
            .O(N__34396),
            .I(N__34312));
    Span4Mux_h I__6615 (
            .O(N__34393),
            .I(N__34301));
    LocalMux I__6614 (
            .O(N__34382),
            .I(N__34301));
    Span4Mux_h I__6613 (
            .O(N__34377),
            .I(N__34301));
    Span4Mux_h I__6612 (
            .O(N__34372),
            .I(N__34301));
    Span4Mux_h I__6611 (
            .O(N__34369),
            .I(N__34301));
    Span12Mux_s10_h I__6610 (
            .O(N__34366),
            .I(N__34298));
    LocalMux I__6609 (
            .O(N__34359),
            .I(N__34291));
    LocalMux I__6608 (
            .O(N__34354),
            .I(N__34291));
    LocalMux I__6607 (
            .O(N__34349),
            .I(N__34291));
    Odrv4 I__6606 (
            .O(N__34346),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__6605 (
            .O(N__34335),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__6604 (
            .O(N__34326),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__6603 (
            .O(N__34317),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__6602 (
            .O(N__34312),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__6601 (
            .O(N__34301),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__6600 (
            .O(N__34298),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__6599 (
            .O(N__34291),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    CascadeMux I__6598 (
            .O(N__34274),
            .I(N__34270));
    InMux I__6597 (
            .O(N__34273),
            .I(N__34265));
    InMux I__6596 (
            .O(N__34270),
            .I(N__34265));
    LocalMux I__6595 (
            .O(N__34265),
            .I(N__34262));
    Odrv12 I__6594 (
            .O(N__34262),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    CEMux I__6593 (
            .O(N__34259),
            .I(N__34255));
    CEMux I__6592 (
            .O(N__34258),
            .I(N__34239));
    LocalMux I__6591 (
            .O(N__34255),
            .I(N__34236));
    InMux I__6590 (
            .O(N__34254),
            .I(N__34229));
    InMux I__6589 (
            .O(N__34253),
            .I(N__34229));
    InMux I__6588 (
            .O(N__34252),
            .I(N__34229));
    CEMux I__6587 (
            .O(N__34251),
            .I(N__34226));
    CEMux I__6586 (
            .O(N__34250),
            .I(N__34223));
    InMux I__6585 (
            .O(N__34249),
            .I(N__34214));
    InMux I__6584 (
            .O(N__34248),
            .I(N__34214));
    InMux I__6583 (
            .O(N__34247),
            .I(N__34214));
    InMux I__6582 (
            .O(N__34246),
            .I(N__34214));
    CEMux I__6581 (
            .O(N__34245),
            .I(N__34211));
    CEMux I__6580 (
            .O(N__34244),
            .I(N__34208));
    CEMux I__6579 (
            .O(N__34243),
            .I(N__34196));
    CEMux I__6578 (
            .O(N__34242),
            .I(N__34193));
    LocalMux I__6577 (
            .O(N__34239),
            .I(N__34186));
    Span4Mux_h I__6576 (
            .O(N__34236),
            .I(N__34170));
    LocalMux I__6575 (
            .O(N__34229),
            .I(N__34170));
    LocalMux I__6574 (
            .O(N__34226),
            .I(N__34167));
    LocalMux I__6573 (
            .O(N__34223),
            .I(N__34156));
    LocalMux I__6572 (
            .O(N__34214),
            .I(N__34156));
    LocalMux I__6571 (
            .O(N__34211),
            .I(N__34156));
    LocalMux I__6570 (
            .O(N__34208),
            .I(N__34152));
    InMux I__6569 (
            .O(N__34207),
            .I(N__34145));
    InMux I__6568 (
            .O(N__34206),
            .I(N__34145));
    InMux I__6567 (
            .O(N__34205),
            .I(N__34145));
    InMux I__6566 (
            .O(N__34204),
            .I(N__34134));
    InMux I__6565 (
            .O(N__34203),
            .I(N__34134));
    InMux I__6564 (
            .O(N__34202),
            .I(N__34134));
    InMux I__6563 (
            .O(N__34201),
            .I(N__34134));
    InMux I__6562 (
            .O(N__34200),
            .I(N__34134));
    CEMux I__6561 (
            .O(N__34199),
            .I(N__34131));
    LocalMux I__6560 (
            .O(N__34196),
            .I(N__34128));
    LocalMux I__6559 (
            .O(N__34193),
            .I(N__34125));
    InMux I__6558 (
            .O(N__34192),
            .I(N__34116));
    InMux I__6557 (
            .O(N__34191),
            .I(N__34116));
    InMux I__6556 (
            .O(N__34190),
            .I(N__34116));
    InMux I__6555 (
            .O(N__34189),
            .I(N__34116));
    Span4Mux_v I__6554 (
            .O(N__34186),
            .I(N__34113));
    CEMux I__6553 (
            .O(N__34185),
            .I(N__34110));
    CEMux I__6552 (
            .O(N__34184),
            .I(N__34107));
    CEMux I__6551 (
            .O(N__34183),
            .I(N__34104));
    InMux I__6550 (
            .O(N__34182),
            .I(N__34095));
    InMux I__6549 (
            .O(N__34181),
            .I(N__34095));
    InMux I__6548 (
            .O(N__34180),
            .I(N__34095));
    InMux I__6547 (
            .O(N__34179),
            .I(N__34095));
    InMux I__6546 (
            .O(N__34178),
            .I(N__34086));
    InMux I__6545 (
            .O(N__34177),
            .I(N__34086));
    InMux I__6544 (
            .O(N__34176),
            .I(N__34086));
    InMux I__6543 (
            .O(N__34175),
            .I(N__34086));
    Span4Mux_v I__6542 (
            .O(N__34170),
            .I(N__34081));
    Span4Mux_v I__6541 (
            .O(N__34167),
            .I(N__34081));
    InMux I__6540 (
            .O(N__34166),
            .I(N__34072));
    InMux I__6539 (
            .O(N__34165),
            .I(N__34072));
    InMux I__6538 (
            .O(N__34164),
            .I(N__34072));
    InMux I__6537 (
            .O(N__34163),
            .I(N__34072));
    Span4Mux_v I__6536 (
            .O(N__34156),
            .I(N__34069));
    CEMux I__6535 (
            .O(N__34155),
            .I(N__34066));
    Span4Mux_h I__6534 (
            .O(N__34152),
            .I(N__34063));
    LocalMux I__6533 (
            .O(N__34145),
            .I(N__34058));
    LocalMux I__6532 (
            .O(N__34134),
            .I(N__34058));
    LocalMux I__6531 (
            .O(N__34131),
            .I(N__34055));
    Span4Mux_h I__6530 (
            .O(N__34128),
            .I(N__34052));
    Span4Mux_v I__6529 (
            .O(N__34125),
            .I(N__34049));
    LocalMux I__6528 (
            .O(N__34116),
            .I(N__34046));
    Span4Mux_v I__6527 (
            .O(N__34113),
            .I(N__34039));
    LocalMux I__6526 (
            .O(N__34110),
            .I(N__34039));
    LocalMux I__6525 (
            .O(N__34107),
            .I(N__34039));
    LocalMux I__6524 (
            .O(N__34104),
            .I(N__34032));
    LocalMux I__6523 (
            .O(N__34095),
            .I(N__34032));
    LocalMux I__6522 (
            .O(N__34086),
            .I(N__34032));
    Span4Mux_h I__6521 (
            .O(N__34081),
            .I(N__34025));
    LocalMux I__6520 (
            .O(N__34072),
            .I(N__34025));
    Span4Mux_h I__6519 (
            .O(N__34069),
            .I(N__34025));
    LocalMux I__6518 (
            .O(N__34066),
            .I(N__34018));
    Span4Mux_h I__6517 (
            .O(N__34063),
            .I(N__34018));
    Span4Mux_h I__6516 (
            .O(N__34058),
            .I(N__34018));
    Span4Mux_h I__6515 (
            .O(N__34055),
            .I(N__34009));
    Span4Mux_h I__6514 (
            .O(N__34052),
            .I(N__34009));
    Span4Mux_h I__6513 (
            .O(N__34049),
            .I(N__34009));
    Span4Mux_h I__6512 (
            .O(N__34046),
            .I(N__34009));
    Span4Mux_v I__6511 (
            .O(N__34039),
            .I(N__34006));
    Span4Mux_v I__6510 (
            .O(N__34032),
            .I(N__34001));
    Span4Mux_v I__6509 (
            .O(N__34025),
            .I(N__34001));
    Span4Mux_v I__6508 (
            .O(N__34018),
            .I(N__33998));
    Span4Mux_v I__6507 (
            .O(N__34009),
            .I(N__33995));
    Odrv4 I__6506 (
            .O(N__34006),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6505 (
            .O(N__34001),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6504 (
            .O(N__33998),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6503 (
            .O(N__33995),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__6502 (
            .O(N__33986),
            .I(N__33983));
    LocalMux I__6501 (
            .O(N__33983),
            .I(N__33979));
    InMux I__6500 (
            .O(N__33982),
            .I(N__33976));
    Odrv4 I__6499 (
            .O(N__33979),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__6498 (
            .O(N__33976),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__6497 (
            .O(N__33971),
            .I(N__33968));
    LocalMux I__6496 (
            .O(N__33968),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__6495 (
            .O(N__33965),
            .I(N__33961));
    InMux I__6494 (
            .O(N__33964),
            .I(N__33958));
    LocalMux I__6493 (
            .O(N__33961),
            .I(N__33955));
    LocalMux I__6492 (
            .O(N__33958),
            .I(N__33952));
    Span4Mux_v I__6491 (
            .O(N__33955),
            .I(N__33948));
    Span4Mux_h I__6490 (
            .O(N__33952),
            .I(N__33945));
    InMux I__6489 (
            .O(N__33951),
            .I(N__33942));
    Odrv4 I__6488 (
            .O(N__33948),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv4 I__6487 (
            .O(N__33945),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    LocalMux I__6486 (
            .O(N__33942),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__6485 (
            .O(N__33935),
            .I(N__33932));
    LocalMux I__6484 (
            .O(N__33932),
            .I(N__33929));
    Span4Mux_v I__6483 (
            .O(N__33929),
            .I(N__33926));
    Odrv4 I__6482 (
            .O(N__33926),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ));
    InMux I__6481 (
            .O(N__33923),
            .I(N__33919));
    InMux I__6480 (
            .O(N__33922),
            .I(N__33916));
    LocalMux I__6479 (
            .O(N__33919),
            .I(N__33913));
    LocalMux I__6478 (
            .O(N__33916),
            .I(N__33909));
    Span4Mux_h I__6477 (
            .O(N__33913),
            .I(N__33906));
    InMux I__6476 (
            .O(N__33912),
            .I(N__33903));
    Odrv12 I__6475 (
            .O(N__33909),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv4 I__6474 (
            .O(N__33906),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    LocalMux I__6473 (
            .O(N__33903),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__6472 (
            .O(N__33896),
            .I(N__33893));
    LocalMux I__6471 (
            .O(N__33893),
            .I(N__33890));
    Odrv12 I__6470 (
            .O(N__33890),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ));
    InMux I__6469 (
            .O(N__33887),
            .I(N__33883));
    CascadeMux I__6468 (
            .O(N__33886),
            .I(N__33880));
    LocalMux I__6467 (
            .O(N__33883),
            .I(N__33877));
    InMux I__6466 (
            .O(N__33880),
            .I(N__33874));
    Span4Mux_h I__6465 (
            .O(N__33877),
            .I(N__33871));
    LocalMux I__6464 (
            .O(N__33874),
            .I(N__33868));
    Span4Mux_h I__6463 (
            .O(N__33871),
            .I(N__33864));
    Span4Mux_h I__6462 (
            .O(N__33868),
            .I(N__33861));
    InMux I__6461 (
            .O(N__33867),
            .I(N__33858));
    Odrv4 I__6460 (
            .O(N__33864),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__6459 (
            .O(N__33861),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    LocalMux I__6458 (
            .O(N__33858),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__6457 (
            .O(N__33851),
            .I(N__33848));
    LocalMux I__6456 (
            .O(N__33848),
            .I(N__33845));
    Odrv12 I__6455 (
            .O(N__33845),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ));
    InMux I__6454 (
            .O(N__33842),
            .I(N__33839));
    LocalMux I__6453 (
            .O(N__33839),
            .I(N__33835));
    InMux I__6452 (
            .O(N__33838),
            .I(N__33832));
    Span4Mux_v I__6451 (
            .O(N__33835),
            .I(N__33829));
    LocalMux I__6450 (
            .O(N__33832),
            .I(N__33826));
    Span4Mux_h I__6449 (
            .O(N__33829),
            .I(N__33820));
    Span4Mux_v I__6448 (
            .O(N__33826),
            .I(N__33820));
    InMux I__6447 (
            .O(N__33825),
            .I(N__33817));
    Odrv4 I__6446 (
            .O(N__33820),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    LocalMux I__6445 (
            .O(N__33817),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__6444 (
            .O(N__33812),
            .I(N__33809));
    LocalMux I__6443 (
            .O(N__33809),
            .I(N__33806));
    Odrv4 I__6442 (
            .O(N__33806),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ));
    InMux I__6441 (
            .O(N__33803),
            .I(N__33800));
    LocalMux I__6440 (
            .O(N__33800),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__6439 (
            .O(N__33797),
            .I(N__33794));
    LocalMux I__6438 (
            .O(N__33794),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__6437 (
            .O(N__33791),
            .I(N__33788));
    LocalMux I__6436 (
            .O(N__33788),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__6435 (
            .O(N__33785),
            .I(N__33782));
    LocalMux I__6434 (
            .O(N__33782),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__6433 (
            .O(N__33779),
            .I(N__33776));
    LocalMux I__6432 (
            .O(N__33776),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__6431 (
            .O(N__33773),
            .I(N__33770));
    LocalMux I__6430 (
            .O(N__33770),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__6429 (
            .O(N__33767),
            .I(N__33764));
    LocalMux I__6428 (
            .O(N__33764),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__6427 (
            .O(N__33761),
            .I(N__33758));
    LocalMux I__6426 (
            .O(N__33758),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__6425 (
            .O(N__33755),
            .I(N__33752));
    LocalMux I__6424 (
            .O(N__33752),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__6423 (
            .O(N__33749),
            .I(N__33746));
    LocalMux I__6422 (
            .O(N__33746),
            .I(N__33743));
    Span4Mux_h I__6421 (
            .O(N__33743),
            .I(N__33740));
    Sp12to4 I__6420 (
            .O(N__33740),
            .I(N__33737));
    Span12Mux_v I__6419 (
            .O(N__33737),
            .I(N__33734));
    Odrv12 I__6418 (
            .O(N__33734),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__6417 (
            .O(N__33731),
            .I(N__33728));
    LocalMux I__6416 (
            .O(N__33728),
            .I(\current_shift_inst.control_input_axb_0 ));
    CascadeMux I__6415 (
            .O(N__33725),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    InMux I__6414 (
            .O(N__33722),
            .I(N__33719));
    LocalMux I__6413 (
            .O(N__33719),
            .I(N__33716));
    Span4Mux_h I__6412 (
            .O(N__33716),
            .I(N__33712));
    InMux I__6411 (
            .O(N__33715),
            .I(N__33709));
    Span4Mux_h I__6410 (
            .O(N__33712),
            .I(N__33706));
    LocalMux I__6409 (
            .O(N__33709),
            .I(N__33703));
    Span4Mux_v I__6408 (
            .O(N__33706),
            .I(N__33700));
    Span4Mux_v I__6407 (
            .O(N__33703),
            .I(N__33697));
    Odrv4 I__6406 (
            .O(N__33700),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv4 I__6405 (
            .O(N__33697),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    CascadeMux I__6404 (
            .O(N__33692),
            .I(N__33687));
    InMux I__6403 (
            .O(N__33691),
            .I(N__33684));
    InMux I__6402 (
            .O(N__33690),
            .I(N__33681));
    InMux I__6401 (
            .O(N__33687),
            .I(N__33678));
    LocalMux I__6400 (
            .O(N__33684),
            .I(\current_shift_inst.N_1326_i ));
    LocalMux I__6399 (
            .O(N__33681),
            .I(\current_shift_inst.N_1326_i ));
    LocalMux I__6398 (
            .O(N__33678),
            .I(\current_shift_inst.N_1326_i ));
    InMux I__6397 (
            .O(N__33671),
            .I(N__33668));
    LocalMux I__6396 (
            .O(N__33668),
            .I(N__33665));
    Odrv4 I__6395 (
            .O(N__33665),
            .I(\current_shift_inst.control_input_axb_12 ));
    CascadeMux I__6394 (
            .O(N__33662),
            .I(\phase_controller_inst1.N_55_cascade_ ));
    InMux I__6393 (
            .O(N__33659),
            .I(N__33656));
    LocalMux I__6392 (
            .O(N__33656),
            .I(N__33653));
    Span4Mux_h I__6391 (
            .O(N__33653),
            .I(N__33649));
    InMux I__6390 (
            .O(N__33652),
            .I(N__33646));
    Odrv4 I__6389 (
            .O(N__33649),
            .I(state_ns_i_a2_1));
    LocalMux I__6388 (
            .O(N__33646),
            .I(state_ns_i_a2_1));
    InMux I__6387 (
            .O(N__33641),
            .I(N__33638));
    LocalMux I__6386 (
            .O(N__33638),
            .I(N__33633));
    InMux I__6385 (
            .O(N__33637),
            .I(N__33630));
    InMux I__6384 (
            .O(N__33636),
            .I(N__33627));
    Span4Mux_v I__6383 (
            .O(N__33633),
            .I(N__33622));
    LocalMux I__6382 (
            .O(N__33630),
            .I(N__33622));
    LocalMux I__6381 (
            .O(N__33627),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    Odrv4 I__6380 (
            .O(N__33622),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    InMux I__6379 (
            .O(N__33617),
            .I(N__33614));
    LocalMux I__6378 (
            .O(N__33614),
            .I(N__33611));
    Span4Mux_v I__6377 (
            .O(N__33611),
            .I(N__33608));
    Span4Mux_h I__6376 (
            .O(N__33608),
            .I(N__33605));
    Odrv4 I__6375 (
            .O(N__33605),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    InMux I__6374 (
            .O(N__33602),
            .I(N__33599));
    LocalMux I__6373 (
            .O(N__33599),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    IoInMux I__6372 (
            .O(N__33596),
            .I(N__33593));
    LocalMux I__6371 (
            .O(N__33593),
            .I(N__33590));
    Span4Mux_s2_v I__6370 (
            .O(N__33590),
            .I(N__33587));
    Sp12to4 I__6369 (
            .O(N__33587),
            .I(N__33584));
    Span12Mux_h I__6368 (
            .O(N__33584),
            .I(N__33580));
    InMux I__6367 (
            .O(N__33583),
            .I(N__33577));
    Odrv12 I__6366 (
            .O(N__33580),
            .I(T23_c));
    LocalMux I__6365 (
            .O(N__33577),
            .I(T23_c));
    InMux I__6364 (
            .O(N__33572),
            .I(N__33566));
    InMux I__6363 (
            .O(N__33571),
            .I(N__33566));
    LocalMux I__6362 (
            .O(N__33566),
            .I(N__33561));
    InMux I__6361 (
            .O(N__33565),
            .I(N__33556));
    InMux I__6360 (
            .O(N__33564),
            .I(N__33556));
    Odrv12 I__6359 (
            .O(N__33561),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__6358 (
            .O(N__33556),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    IoInMux I__6357 (
            .O(N__33551),
            .I(N__33548));
    LocalMux I__6356 (
            .O(N__33548),
            .I(N__33545));
    IoSpan4Mux I__6355 (
            .O(N__33545),
            .I(N__33542));
    Span4Mux_s3_v I__6354 (
            .O(N__33542),
            .I(N__33539));
    Span4Mux_v I__6353 (
            .O(N__33539),
            .I(N__33536));
    Span4Mux_v I__6352 (
            .O(N__33536),
            .I(N__33532));
    InMux I__6351 (
            .O(N__33535),
            .I(N__33529));
    Odrv4 I__6350 (
            .O(N__33532),
            .I(T45_c));
    LocalMux I__6349 (
            .O(N__33529),
            .I(T45_c));
    InMux I__6348 (
            .O(N__33524),
            .I(N__33520));
    InMux I__6347 (
            .O(N__33523),
            .I(N__33517));
    LocalMux I__6346 (
            .O(N__33520),
            .I(N__33514));
    LocalMux I__6345 (
            .O(N__33517),
            .I(N__33511));
    Span4Mux_h I__6344 (
            .O(N__33514),
            .I(N__33508));
    Span12Mux_v I__6343 (
            .O(N__33511),
            .I(N__33504));
    Span4Mux_v I__6342 (
            .O(N__33508),
            .I(N__33501));
    InMux I__6341 (
            .O(N__33507),
            .I(N__33498));
    Odrv12 I__6340 (
            .O(N__33504),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__6339 (
            .O(N__33501),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    LocalMux I__6338 (
            .O(N__33498),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__6337 (
            .O(N__33491),
            .I(N__33488));
    LocalMux I__6336 (
            .O(N__33488),
            .I(N__33485));
    Odrv4 I__6335 (
            .O(N__33485),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ));
    CascadeMux I__6334 (
            .O(N__33482),
            .I(N__33478));
    InMux I__6333 (
            .O(N__33481),
            .I(N__33475));
    InMux I__6332 (
            .O(N__33478),
            .I(N__33472));
    LocalMux I__6331 (
            .O(N__33475),
            .I(N__33469));
    LocalMux I__6330 (
            .O(N__33472),
            .I(N__33466));
    Span4Mux_v I__6329 (
            .O(N__33469),
            .I(N__33462));
    Span4Mux_h I__6328 (
            .O(N__33466),
            .I(N__33459));
    InMux I__6327 (
            .O(N__33465),
            .I(N__33456));
    Odrv4 I__6326 (
            .O(N__33462),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__6325 (
            .O(N__33459),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    LocalMux I__6324 (
            .O(N__33456),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__6323 (
            .O(N__33449),
            .I(N__33446));
    LocalMux I__6322 (
            .O(N__33446),
            .I(N__33443));
    Odrv4 I__6321 (
            .O(N__33443),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ));
    InMux I__6320 (
            .O(N__33440),
            .I(N__33436));
    InMux I__6319 (
            .O(N__33439),
            .I(N__33433));
    LocalMux I__6318 (
            .O(N__33436),
            .I(N__33427));
    LocalMux I__6317 (
            .O(N__33433),
            .I(N__33427));
    InMux I__6316 (
            .O(N__33432),
            .I(N__33424));
    Span4Mux_h I__6315 (
            .O(N__33427),
            .I(N__33421));
    LocalMux I__6314 (
            .O(N__33424),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv4 I__6313 (
            .O(N__33421),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    CascadeMux I__6312 (
            .O(N__33416),
            .I(N__33413));
    InMux I__6311 (
            .O(N__33413),
            .I(N__33409));
    InMux I__6310 (
            .O(N__33412),
            .I(N__33406));
    LocalMux I__6309 (
            .O(N__33409),
            .I(N__33400));
    LocalMux I__6308 (
            .O(N__33406),
            .I(N__33400));
    InMux I__6307 (
            .O(N__33405),
            .I(N__33397));
    Span4Mux_h I__6306 (
            .O(N__33400),
            .I(N__33394));
    LocalMux I__6305 (
            .O(N__33397),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    Odrv4 I__6304 (
            .O(N__33394),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    InMux I__6303 (
            .O(N__33389),
            .I(N__33385));
    InMux I__6302 (
            .O(N__33388),
            .I(N__33382));
    LocalMux I__6301 (
            .O(N__33385),
            .I(N__33379));
    LocalMux I__6300 (
            .O(N__33382),
            .I(N__33376));
    Span4Mux_v I__6299 (
            .O(N__33379),
            .I(N__33373));
    Span4Mux_h I__6298 (
            .O(N__33376),
            .I(N__33369));
    Span4Mux_h I__6297 (
            .O(N__33373),
            .I(N__33366));
    InMux I__6296 (
            .O(N__33372),
            .I(N__33363));
    Odrv4 I__6295 (
            .O(N__33369),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__6294 (
            .O(N__33366),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    LocalMux I__6293 (
            .O(N__33363),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__6292 (
            .O(N__33356),
            .I(N__33353));
    LocalMux I__6291 (
            .O(N__33353),
            .I(N__33350));
    Odrv4 I__6290 (
            .O(N__33350),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ));
    InMux I__6289 (
            .O(N__33347),
            .I(N__33344));
    LocalMux I__6288 (
            .O(N__33344),
            .I(N__33339));
    InMux I__6287 (
            .O(N__33343),
            .I(N__33336));
    InMux I__6286 (
            .O(N__33342),
            .I(N__33333));
    Span4Mux_v I__6285 (
            .O(N__33339),
            .I(N__33328));
    LocalMux I__6284 (
            .O(N__33336),
            .I(N__33328));
    LocalMux I__6283 (
            .O(N__33333),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    Odrv4 I__6282 (
            .O(N__33328),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    InMux I__6281 (
            .O(N__33323),
            .I(N__33320));
    LocalMux I__6280 (
            .O(N__33320),
            .I(N__33315));
    InMux I__6279 (
            .O(N__33319),
            .I(N__33312));
    InMux I__6278 (
            .O(N__33318),
            .I(N__33309));
    Span4Mux_v I__6277 (
            .O(N__33315),
            .I(N__33304));
    LocalMux I__6276 (
            .O(N__33312),
            .I(N__33304));
    LocalMux I__6275 (
            .O(N__33309),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    Odrv4 I__6274 (
            .O(N__33304),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    CascadeMux I__6273 (
            .O(N__33299),
            .I(N__33295));
    InMux I__6272 (
            .O(N__33298),
            .I(N__33292));
    InMux I__6271 (
            .O(N__33295),
            .I(N__33289));
    LocalMux I__6270 (
            .O(N__33292),
            .I(N__33286));
    LocalMux I__6269 (
            .O(N__33289),
            .I(N__33283));
    Span4Mux_h I__6268 (
            .O(N__33286),
            .I(N__33279));
    Span4Mux_v I__6267 (
            .O(N__33283),
            .I(N__33276));
    InMux I__6266 (
            .O(N__33282),
            .I(N__33273));
    Odrv4 I__6265 (
            .O(N__33279),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv4 I__6264 (
            .O(N__33276),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    LocalMux I__6263 (
            .O(N__33273),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__6262 (
            .O(N__33266),
            .I(N__33263));
    LocalMux I__6261 (
            .O(N__33263),
            .I(N__33260));
    Odrv4 I__6260 (
            .O(N__33260),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    InMux I__6259 (
            .O(N__33257),
            .I(N__33254));
    LocalMux I__6258 (
            .O(N__33254),
            .I(N__33251));
    Odrv4 I__6257 (
            .O(N__33251),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__6256 (
            .O(N__33248),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__6255 (
            .O(N__33245),
            .I(N__33242));
    LocalMux I__6254 (
            .O(N__33242),
            .I(N__33239));
    Odrv4 I__6253 (
            .O(N__33239),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__6252 (
            .O(N__33236),
            .I(bfn_12_14_0_));
    InMux I__6251 (
            .O(N__33233),
            .I(N__33230));
    LocalMux I__6250 (
            .O(N__33230),
            .I(N__33227));
    Odrv12 I__6249 (
            .O(N__33227),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__6248 (
            .O(N__33224),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__6247 (
            .O(N__33221),
            .I(N__33218));
    LocalMux I__6246 (
            .O(N__33218),
            .I(N__33215));
    Odrv4 I__6245 (
            .O(N__33215),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__6244 (
            .O(N__33212),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__6243 (
            .O(N__33209),
            .I(N__33206));
    LocalMux I__6242 (
            .O(N__33206),
            .I(N__33203));
    Odrv4 I__6241 (
            .O(N__33203),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__6240 (
            .O(N__33200),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__6239 (
            .O(N__33197),
            .I(N__33194));
    LocalMux I__6238 (
            .O(N__33194),
            .I(N__33191));
    Odrv12 I__6237 (
            .O(N__33191),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__6236 (
            .O(N__33188),
            .I(N__33181));
    InMux I__6235 (
            .O(N__33187),
            .I(N__33181));
    InMux I__6234 (
            .O(N__33186),
            .I(N__33178));
    LocalMux I__6233 (
            .O(N__33181),
            .I(N__33175));
    LocalMux I__6232 (
            .O(N__33178),
            .I(N__33172));
    Span4Mux_h I__6231 (
            .O(N__33175),
            .I(N__33169));
    Odrv12 I__6230 (
            .O(N__33172),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__6229 (
            .O(N__33169),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__6228 (
            .O(N__33164),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__6227 (
            .O(N__33161),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__6226 (
            .O(N__33158),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__6225 (
            .O(N__33155),
            .I(N__33152));
    LocalMux I__6224 (
            .O(N__33152),
            .I(N__33148));
    InMux I__6223 (
            .O(N__33151),
            .I(N__33145));
    Span4Mux_h I__6222 (
            .O(N__33148),
            .I(N__33142));
    LocalMux I__6221 (
            .O(N__33145),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv4 I__6220 (
            .O(N__33142),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__6219 (
            .O(N__33137),
            .I(N__33134));
    LocalMux I__6218 (
            .O(N__33134),
            .I(N__33131));
    Span4Mux_v I__6217 (
            .O(N__33131),
            .I(N__33128));
    Span4Mux_h I__6216 (
            .O(N__33128),
            .I(N__33125));
    Odrv4 I__6215 (
            .O(N__33125),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__6214 (
            .O(N__33122),
            .I(N__33119));
    LocalMux I__6213 (
            .O(N__33119),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__6212 (
            .O(N__33116),
            .I(N__33113));
    LocalMux I__6211 (
            .O(N__33113),
            .I(N__33110));
    Odrv4 I__6210 (
            .O(N__33110),
            .I(\current_shift_inst.control_input_18 ));
    InMux I__6209 (
            .O(N__33107),
            .I(N__33104));
    LocalMux I__6208 (
            .O(N__33104),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__6207 (
            .O(N__33101),
            .I(N__33098));
    LocalMux I__6206 (
            .O(N__33098),
            .I(N__33095));
    Odrv4 I__6205 (
            .O(N__33095),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__6204 (
            .O(N__33092),
            .I(N__33089));
    LocalMux I__6203 (
            .O(N__33089),
            .I(N__33085));
    InMux I__6202 (
            .O(N__33088),
            .I(N__33082));
    Span4Mux_h I__6201 (
            .O(N__33085),
            .I(N__33077));
    LocalMux I__6200 (
            .O(N__33082),
            .I(N__33077));
    Span4Mux_h I__6199 (
            .O(N__33077),
            .I(N__33074));
    Odrv4 I__6198 (
            .O(N__33074),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__6197 (
            .O(N__33071),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    CascadeMux I__6196 (
            .O(N__33068),
            .I(N__33065));
    InMux I__6195 (
            .O(N__33065),
            .I(N__33062));
    LocalMux I__6194 (
            .O(N__33062),
            .I(N__33059));
    Odrv4 I__6193 (
            .O(N__33059),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__6192 (
            .O(N__33056),
            .I(N__33053));
    LocalMux I__6191 (
            .O(N__33053),
            .I(N__33049));
    InMux I__6190 (
            .O(N__33052),
            .I(N__33046));
    Span4Mux_h I__6189 (
            .O(N__33049),
            .I(N__33041));
    LocalMux I__6188 (
            .O(N__33046),
            .I(N__33041));
    Span4Mux_h I__6187 (
            .O(N__33041),
            .I(N__33038));
    Odrv4 I__6186 (
            .O(N__33038),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__6185 (
            .O(N__33035),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__6184 (
            .O(N__33032),
            .I(N__33029));
    LocalMux I__6183 (
            .O(N__33029),
            .I(N__33026));
    Odrv4 I__6182 (
            .O(N__33026),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__6181 (
            .O(N__33023),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__6180 (
            .O(N__33020),
            .I(N__33017));
    LocalMux I__6179 (
            .O(N__33017),
            .I(N__33014));
    Odrv12 I__6178 (
            .O(N__33014),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__6177 (
            .O(N__33011),
            .I(N__33008));
    LocalMux I__6176 (
            .O(N__33008),
            .I(N__33003));
    InMux I__6175 (
            .O(N__33007),
            .I(N__32998));
    InMux I__6174 (
            .O(N__33006),
            .I(N__32998));
    Span4Mux_v I__6173 (
            .O(N__33003),
            .I(N__32995));
    LocalMux I__6172 (
            .O(N__32998),
            .I(N__32992));
    Span4Mux_h I__6171 (
            .O(N__32995),
            .I(N__32987));
    Span4Mux_v I__6170 (
            .O(N__32992),
            .I(N__32987));
    Odrv4 I__6169 (
            .O(N__32987),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__6168 (
            .O(N__32984),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__6167 (
            .O(N__32981),
            .I(N__32978));
    LocalMux I__6166 (
            .O(N__32978),
            .I(N__32975));
    Odrv4 I__6165 (
            .O(N__32975),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__6164 (
            .O(N__32972),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__6163 (
            .O(N__32969),
            .I(N__32966));
    LocalMux I__6162 (
            .O(N__32966),
            .I(N__32963));
    Odrv4 I__6161 (
            .O(N__32963),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__6160 (
            .O(N__32960),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__6159 (
            .O(N__32957),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__6158 (
            .O(N__32954),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__6157 (
            .O(N__32951),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__6156 (
            .O(N__32948),
            .I(bfn_12_12_0_));
    InMux I__6155 (
            .O(N__32945),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__6154 (
            .O(N__32942),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__6153 (
            .O(N__32939),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__6152 (
            .O(N__32936),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__6151 (
            .O(N__32933),
            .I(\current_shift_inst.control_input_cry_12 ));
    CascadeMux I__6150 (
            .O(N__32930),
            .I(N__32926));
    InMux I__6149 (
            .O(N__32929),
            .I(N__32923));
    InMux I__6148 (
            .O(N__32926),
            .I(N__32918));
    LocalMux I__6147 (
            .O(N__32923),
            .I(N__32915));
    CascadeMux I__6146 (
            .O(N__32922),
            .I(N__32912));
    InMux I__6145 (
            .O(N__32921),
            .I(N__32909));
    LocalMux I__6144 (
            .O(N__32918),
            .I(N__32906));
    Span4Mux_h I__6143 (
            .O(N__32915),
            .I(N__32903));
    InMux I__6142 (
            .O(N__32912),
            .I(N__32900));
    LocalMux I__6141 (
            .O(N__32909),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv12 I__6140 (
            .O(N__32906),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv4 I__6139 (
            .O(N__32903),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__6138 (
            .O(N__32900),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__6137 (
            .O(N__32891),
            .I(N__32888));
    LocalMux I__6136 (
            .O(N__32888),
            .I(N__32884));
    InMux I__6135 (
            .O(N__32887),
            .I(N__32880));
    Span4Mux_h I__6134 (
            .O(N__32884),
            .I(N__32877));
    InMux I__6133 (
            .O(N__32883),
            .I(N__32874));
    LocalMux I__6132 (
            .O(N__32880),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    Odrv4 I__6131 (
            .O(N__32877),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    LocalMux I__6130 (
            .O(N__32874),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    InMux I__6129 (
            .O(N__32867),
            .I(N__32863));
    InMux I__6128 (
            .O(N__32866),
            .I(N__32860));
    LocalMux I__6127 (
            .O(N__32863),
            .I(N__32857));
    LocalMux I__6126 (
            .O(N__32860),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    Odrv12 I__6125 (
            .O(N__32857),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    CascadeMux I__6124 (
            .O(N__32852),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_));
    InMux I__6123 (
            .O(N__32849),
            .I(N__32843));
    InMux I__6122 (
            .O(N__32848),
            .I(N__32843));
    LocalMux I__6121 (
            .O(N__32843),
            .I(N__32839));
    InMux I__6120 (
            .O(N__32842),
            .I(N__32835));
    Span4Mux_h I__6119 (
            .O(N__32839),
            .I(N__32832));
    InMux I__6118 (
            .O(N__32838),
            .I(N__32829));
    LocalMux I__6117 (
            .O(N__32835),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    Odrv4 I__6116 (
            .O(N__32832),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    LocalMux I__6115 (
            .O(N__32829),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__6114 (
            .O(N__32822),
            .I(N__32819));
    LocalMux I__6113 (
            .O(N__32819),
            .I(N__32816));
    Span4Mux_v I__6112 (
            .O(N__32816),
            .I(N__32813));
    Odrv4 I__6111 (
            .O(N__32813),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__6110 (
            .O(N__32810),
            .I(N__32806));
    InMux I__6109 (
            .O(N__32809),
            .I(N__32801));
    LocalMux I__6108 (
            .O(N__32806),
            .I(N__32798));
    CascadeMux I__6107 (
            .O(N__32805),
            .I(N__32795));
    InMux I__6106 (
            .O(N__32804),
            .I(N__32792));
    LocalMux I__6105 (
            .O(N__32801),
            .I(N__32787));
    Span4Mux_v I__6104 (
            .O(N__32798),
            .I(N__32787));
    InMux I__6103 (
            .O(N__32795),
            .I(N__32784));
    LocalMux I__6102 (
            .O(N__32792),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv4 I__6101 (
            .O(N__32787),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__6100 (
            .O(N__32784),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__6099 (
            .O(N__32777),
            .I(N__32774));
    LocalMux I__6098 (
            .O(N__32774),
            .I(N__32770));
    InMux I__6097 (
            .O(N__32773),
            .I(N__32766));
    Span4Mux_h I__6096 (
            .O(N__32770),
            .I(N__32763));
    InMux I__6095 (
            .O(N__32769),
            .I(N__32760));
    LocalMux I__6094 (
            .O(N__32766),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    Odrv4 I__6093 (
            .O(N__32763),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    LocalMux I__6092 (
            .O(N__32760),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    InMux I__6091 (
            .O(N__32753),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__6090 (
            .O(N__32750),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__6089 (
            .O(N__32747),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__6088 (
            .O(N__32744),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__6087 (
            .O(N__32741),
            .I(N__32738));
    LocalMux I__6086 (
            .O(N__32738),
            .I(il_min_comp1_D1));
    InMux I__6085 (
            .O(N__32735),
            .I(N__32732));
    LocalMux I__6084 (
            .O(N__32732),
            .I(N__32727));
    InMux I__6083 (
            .O(N__32731),
            .I(N__32724));
    InMux I__6082 (
            .O(N__32730),
            .I(N__32721));
    Span4Mux_v I__6081 (
            .O(N__32727),
            .I(N__32718));
    LocalMux I__6080 (
            .O(N__32724),
            .I(N__32713));
    LocalMux I__6079 (
            .O(N__32721),
            .I(N__32713));
    Odrv4 I__6078 (
            .O(N__32718),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    Odrv12 I__6077 (
            .O(N__32713),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    InMux I__6076 (
            .O(N__32708),
            .I(N__32704));
    InMux I__6075 (
            .O(N__32707),
            .I(N__32701));
    LocalMux I__6074 (
            .O(N__32704),
            .I(N__32696));
    LocalMux I__6073 (
            .O(N__32701),
            .I(N__32693));
    CascadeMux I__6072 (
            .O(N__32700),
            .I(N__32690));
    InMux I__6071 (
            .O(N__32699),
            .I(N__32687));
    Span4Mux_h I__6070 (
            .O(N__32696),
            .I(N__32682));
    Span4Mux_h I__6069 (
            .O(N__32693),
            .I(N__32682));
    InMux I__6068 (
            .O(N__32690),
            .I(N__32679));
    LocalMux I__6067 (
            .O(N__32687),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv4 I__6066 (
            .O(N__32682),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    LocalMux I__6065 (
            .O(N__32679),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__6064 (
            .O(N__32672),
            .I(N__32666));
    InMux I__6063 (
            .O(N__32671),
            .I(N__32666));
    LocalMux I__6062 (
            .O(N__32666),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ));
    InMux I__6061 (
            .O(N__32663),
            .I(N__32659));
    InMux I__6060 (
            .O(N__32662),
            .I(N__32655));
    LocalMux I__6059 (
            .O(N__32659),
            .I(N__32652));
    InMux I__6058 (
            .O(N__32658),
            .I(N__32649));
    LocalMux I__6057 (
            .O(N__32655),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    Odrv12 I__6056 (
            .O(N__32652),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__6055 (
            .O(N__32649),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    InMux I__6054 (
            .O(N__32642),
            .I(N__32639));
    LocalMux I__6053 (
            .O(N__32639),
            .I(N__32635));
    InMux I__6052 (
            .O(N__32638),
            .I(N__32631));
    Span4Mux_h I__6051 (
            .O(N__32635),
            .I(N__32627));
    InMux I__6050 (
            .O(N__32634),
            .I(N__32624));
    LocalMux I__6049 (
            .O(N__32631),
            .I(N__32621));
    InMux I__6048 (
            .O(N__32630),
            .I(N__32618));
    Odrv4 I__6047 (
            .O(N__32627),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__6046 (
            .O(N__32624),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    Odrv12 I__6045 (
            .O(N__32621),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__6044 (
            .O(N__32618),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__6043 (
            .O(N__32609),
            .I(N__32606));
    LocalMux I__6042 (
            .O(N__32606),
            .I(N__32603));
    Span4Mux_v I__6041 (
            .O(N__32603),
            .I(N__32600));
    Odrv4 I__6040 (
            .O(N__32600),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    InMux I__6039 (
            .O(N__32597),
            .I(N__32594));
    LocalMux I__6038 (
            .O(N__32594),
            .I(N__32591));
    Span4Mux_v I__6037 (
            .O(N__32591),
            .I(N__32588));
    Odrv4 I__6036 (
            .O(N__32588),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    CascadeMux I__6035 (
            .O(N__32585),
            .I(N__32581));
    InMux I__6034 (
            .O(N__32584),
            .I(N__32577));
    InMux I__6033 (
            .O(N__32581),
            .I(N__32574));
    InMux I__6032 (
            .O(N__32580),
            .I(N__32571));
    LocalMux I__6031 (
            .O(N__32577),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__6030 (
            .O(N__32574),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__6029 (
            .O(N__32571),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__6028 (
            .O(N__32564),
            .I(N__32559));
    InMux I__6027 (
            .O(N__32563),
            .I(N__32554));
    InMux I__6026 (
            .O(N__32562),
            .I(N__32554));
    LocalMux I__6025 (
            .O(N__32559),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__6024 (
            .O(N__32554),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__6023 (
            .O(N__32549),
            .I(N__32545));
    InMux I__6022 (
            .O(N__32548),
            .I(N__32540));
    InMux I__6021 (
            .O(N__32545),
            .I(N__32540));
    LocalMux I__6020 (
            .O(N__32540),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__6019 (
            .O(N__32537),
            .I(N__32533));
    InMux I__6018 (
            .O(N__32536),
            .I(N__32530));
    LocalMux I__6017 (
            .O(N__32533),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    LocalMux I__6016 (
            .O(N__32530),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__6015 (
            .O(N__32525),
            .I(N__32522));
    InMux I__6014 (
            .O(N__32522),
            .I(N__32519));
    LocalMux I__6013 (
            .O(N__32519),
            .I(N__32516));
    Span4Mux_v I__6012 (
            .O(N__32516),
            .I(N__32513));
    Span4Mux_h I__6011 (
            .O(N__32513),
            .I(N__32510));
    Odrv4 I__6010 (
            .O(N__32510),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    InMux I__6009 (
            .O(N__32507),
            .I(N__32504));
    LocalMux I__6008 (
            .O(N__32504),
            .I(N__32500));
    InMux I__6007 (
            .O(N__32503),
            .I(N__32496));
    Span4Mux_h I__6006 (
            .O(N__32500),
            .I(N__32493));
    InMux I__6005 (
            .O(N__32499),
            .I(N__32490));
    LocalMux I__6004 (
            .O(N__32496),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv4 I__6003 (
            .O(N__32493),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    LocalMux I__6002 (
            .O(N__32490),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    InMux I__6001 (
            .O(N__32483),
            .I(N__32480));
    LocalMux I__6000 (
            .O(N__32480),
            .I(N__32476));
    InMux I__5999 (
            .O(N__32479),
            .I(N__32472));
    Span4Mux_v I__5998 (
            .O(N__32476),
            .I(N__32469));
    InMux I__5997 (
            .O(N__32475),
            .I(N__32466));
    LocalMux I__5996 (
            .O(N__32472),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    Odrv4 I__5995 (
            .O(N__32469),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    LocalMux I__5994 (
            .O(N__32466),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    InMux I__5993 (
            .O(N__32459),
            .I(N__32456));
    LocalMux I__5992 (
            .O(N__32456),
            .I(N__32452));
    InMux I__5991 (
            .O(N__32455),
            .I(N__32448));
    Span4Mux_h I__5990 (
            .O(N__32452),
            .I(N__32445));
    InMux I__5989 (
            .O(N__32451),
            .I(N__32442));
    LocalMux I__5988 (
            .O(N__32448),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    Odrv4 I__5987 (
            .O(N__32445),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    LocalMux I__5986 (
            .O(N__32442),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    CascadeMux I__5985 (
            .O(N__32435),
            .I(N__32432));
    InMux I__5984 (
            .O(N__32432),
            .I(N__32429));
    LocalMux I__5983 (
            .O(N__32429),
            .I(N__32425));
    InMux I__5982 (
            .O(N__32428),
            .I(N__32421));
    Span4Mux_h I__5981 (
            .O(N__32425),
            .I(N__32418));
    InMux I__5980 (
            .O(N__32424),
            .I(N__32415));
    LocalMux I__5979 (
            .O(N__32421),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    Odrv4 I__5978 (
            .O(N__32418),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    LocalMux I__5977 (
            .O(N__32415),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    InMux I__5976 (
            .O(N__32408),
            .I(N__32405));
    LocalMux I__5975 (
            .O(N__32405),
            .I(N__32402));
    Odrv4 I__5974 (
            .O(N__32402),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    CascadeMux I__5973 (
            .O(N__32399),
            .I(N__32376));
    CascadeMux I__5972 (
            .O(N__32398),
            .I(N__32373));
    InMux I__5971 (
            .O(N__32397),
            .I(N__32370));
    CascadeMux I__5970 (
            .O(N__32396),
            .I(N__32362));
    CascadeMux I__5969 (
            .O(N__32395),
            .I(N__32359));
    CascadeMux I__5968 (
            .O(N__32394),
            .I(N__32356));
    CascadeMux I__5967 (
            .O(N__32393),
            .I(N__32353));
    InMux I__5966 (
            .O(N__32392),
            .I(N__32343));
    InMux I__5965 (
            .O(N__32391),
            .I(N__32343));
    InMux I__5964 (
            .O(N__32390),
            .I(N__32343));
    InMux I__5963 (
            .O(N__32389),
            .I(N__32332));
    InMux I__5962 (
            .O(N__32388),
            .I(N__32332));
    InMux I__5961 (
            .O(N__32387),
            .I(N__32332));
    InMux I__5960 (
            .O(N__32386),
            .I(N__32332));
    InMux I__5959 (
            .O(N__32385),
            .I(N__32332));
    InMux I__5958 (
            .O(N__32384),
            .I(N__32329));
    CascadeMux I__5957 (
            .O(N__32383),
            .I(N__32323));
    CascadeMux I__5956 (
            .O(N__32382),
            .I(N__32320));
    InMux I__5955 (
            .O(N__32381),
            .I(N__32309));
    InMux I__5954 (
            .O(N__32380),
            .I(N__32309));
    InMux I__5953 (
            .O(N__32379),
            .I(N__32309));
    InMux I__5952 (
            .O(N__32376),
            .I(N__32309));
    InMux I__5951 (
            .O(N__32373),
            .I(N__32309));
    LocalMux I__5950 (
            .O(N__32370),
            .I(N__32306));
    InMux I__5949 (
            .O(N__32369),
            .I(N__32299));
    InMux I__5948 (
            .O(N__32368),
            .I(N__32299));
    InMux I__5947 (
            .O(N__32367),
            .I(N__32299));
    InMux I__5946 (
            .O(N__32366),
            .I(N__32292));
    InMux I__5945 (
            .O(N__32365),
            .I(N__32292));
    InMux I__5944 (
            .O(N__32362),
            .I(N__32292));
    InMux I__5943 (
            .O(N__32359),
            .I(N__32279));
    InMux I__5942 (
            .O(N__32356),
            .I(N__32279));
    InMux I__5941 (
            .O(N__32353),
            .I(N__32279));
    InMux I__5940 (
            .O(N__32352),
            .I(N__32279));
    InMux I__5939 (
            .O(N__32351),
            .I(N__32279));
    InMux I__5938 (
            .O(N__32350),
            .I(N__32279));
    LocalMux I__5937 (
            .O(N__32343),
            .I(N__32276));
    LocalMux I__5936 (
            .O(N__32332),
            .I(N__32273));
    LocalMux I__5935 (
            .O(N__32329),
            .I(N__32270));
    InMux I__5934 (
            .O(N__32328),
            .I(N__32259));
    InMux I__5933 (
            .O(N__32327),
            .I(N__32259));
    InMux I__5932 (
            .O(N__32326),
            .I(N__32259));
    InMux I__5931 (
            .O(N__32323),
            .I(N__32259));
    InMux I__5930 (
            .O(N__32320),
            .I(N__32259));
    LocalMux I__5929 (
            .O(N__32309),
            .I(N__32254));
    Span4Mux_v I__5928 (
            .O(N__32306),
            .I(N__32254));
    LocalMux I__5927 (
            .O(N__32299),
            .I(N__32249));
    LocalMux I__5926 (
            .O(N__32292),
            .I(N__32249));
    LocalMux I__5925 (
            .O(N__32279),
            .I(N__32246));
    Span4Mux_v I__5924 (
            .O(N__32276),
            .I(N__32241));
    Span4Mux_v I__5923 (
            .O(N__32273),
            .I(N__32241));
    Span4Mux_v I__5922 (
            .O(N__32270),
            .I(N__32238));
    LocalMux I__5921 (
            .O(N__32259),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__5920 (
            .O(N__32254),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv12 I__5919 (
            .O(N__32249),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__5918 (
            .O(N__32246),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__5917 (
            .O(N__32241),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__5916 (
            .O(N__32238),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    CascadeMux I__5915 (
            .O(N__32225),
            .I(N__32220));
    CascadeMux I__5914 (
            .O(N__32224),
            .I(N__32216));
    CascadeMux I__5913 (
            .O(N__32223),
            .I(N__32208));
    InMux I__5912 (
            .O(N__32220),
            .I(N__32205));
    CascadeMux I__5911 (
            .O(N__32219),
            .I(N__32194));
    InMux I__5910 (
            .O(N__32216),
            .I(N__32189));
    CascadeMux I__5909 (
            .O(N__32215),
            .I(N__32184));
    CascadeMux I__5908 (
            .O(N__32214),
            .I(N__32181));
    CascadeMux I__5907 (
            .O(N__32213),
            .I(N__32178));
    InMux I__5906 (
            .O(N__32212),
            .I(N__32171));
    InMux I__5905 (
            .O(N__32211),
            .I(N__32171));
    InMux I__5904 (
            .O(N__32208),
            .I(N__32171));
    LocalMux I__5903 (
            .O(N__32205),
            .I(N__32168));
    CascadeMux I__5902 (
            .O(N__32204),
            .I(N__32165));
    CascadeMux I__5901 (
            .O(N__32203),
            .I(N__32162));
    CascadeMux I__5900 (
            .O(N__32202),
            .I(N__32159));
    InMux I__5899 (
            .O(N__32201),
            .I(N__32142));
    InMux I__5898 (
            .O(N__32200),
            .I(N__32142));
    InMux I__5897 (
            .O(N__32199),
            .I(N__32142));
    InMux I__5896 (
            .O(N__32198),
            .I(N__32142));
    InMux I__5895 (
            .O(N__32197),
            .I(N__32142));
    InMux I__5894 (
            .O(N__32194),
            .I(N__32135));
    InMux I__5893 (
            .O(N__32193),
            .I(N__32135));
    InMux I__5892 (
            .O(N__32192),
            .I(N__32135));
    LocalMux I__5891 (
            .O(N__32189),
            .I(N__32127));
    InMux I__5890 (
            .O(N__32188),
            .I(N__32116));
    InMux I__5889 (
            .O(N__32187),
            .I(N__32116));
    InMux I__5888 (
            .O(N__32184),
            .I(N__32116));
    InMux I__5887 (
            .O(N__32181),
            .I(N__32116));
    InMux I__5886 (
            .O(N__32178),
            .I(N__32116));
    LocalMux I__5885 (
            .O(N__32171),
            .I(N__32113));
    Span4Mux_v I__5884 (
            .O(N__32168),
            .I(N__32110));
    InMux I__5883 (
            .O(N__32165),
            .I(N__32103));
    InMux I__5882 (
            .O(N__32162),
            .I(N__32103));
    InMux I__5881 (
            .O(N__32159),
            .I(N__32103));
    InMux I__5880 (
            .O(N__32158),
            .I(N__32096));
    InMux I__5879 (
            .O(N__32157),
            .I(N__32096));
    InMux I__5878 (
            .O(N__32156),
            .I(N__32096));
    InMux I__5877 (
            .O(N__32155),
            .I(N__32089));
    InMux I__5876 (
            .O(N__32154),
            .I(N__32089));
    InMux I__5875 (
            .O(N__32153),
            .I(N__32089));
    LocalMux I__5874 (
            .O(N__32142),
            .I(N__32084));
    LocalMux I__5873 (
            .O(N__32135),
            .I(N__32084));
    InMux I__5872 (
            .O(N__32134),
            .I(N__32073));
    InMux I__5871 (
            .O(N__32133),
            .I(N__32073));
    InMux I__5870 (
            .O(N__32132),
            .I(N__32073));
    InMux I__5869 (
            .O(N__32131),
            .I(N__32073));
    InMux I__5868 (
            .O(N__32130),
            .I(N__32073));
    Sp12to4 I__5867 (
            .O(N__32127),
            .I(N__32068));
    LocalMux I__5866 (
            .O(N__32116),
            .I(N__32068));
    Span4Mux_h I__5865 (
            .O(N__32113),
            .I(N__32065));
    Sp12to4 I__5864 (
            .O(N__32110),
            .I(N__32056));
    LocalMux I__5863 (
            .O(N__32103),
            .I(N__32056));
    LocalMux I__5862 (
            .O(N__32096),
            .I(N__32056));
    LocalMux I__5861 (
            .O(N__32089),
            .I(N__32056));
    Span4Mux_v I__5860 (
            .O(N__32084),
            .I(N__32053));
    LocalMux I__5859 (
            .O(N__32073),
            .I(N__32048));
    Span12Mux_v I__5858 (
            .O(N__32068),
            .I(N__32048));
    Span4Mux_v I__5857 (
            .O(N__32065),
            .I(N__32045));
    Span12Mux_h I__5856 (
            .O(N__32056),
            .I(N__32042));
    Odrv4 I__5855 (
            .O(N__32053),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv12 I__5854 (
            .O(N__32048),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__5853 (
            .O(N__32045),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv12 I__5852 (
            .O(N__32042),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    InMux I__5851 (
            .O(N__32033),
            .I(N__32010));
    InMux I__5850 (
            .O(N__32032),
            .I(N__32006));
    InMux I__5849 (
            .O(N__32031),
            .I(N__32000));
    InMux I__5848 (
            .O(N__32030),
            .I(N__31993));
    InMux I__5847 (
            .O(N__32029),
            .I(N__31993));
    InMux I__5846 (
            .O(N__32028),
            .I(N__31993));
    InMux I__5845 (
            .O(N__32027),
            .I(N__31981));
    InMux I__5844 (
            .O(N__32026),
            .I(N__31981));
    InMux I__5843 (
            .O(N__32025),
            .I(N__31981));
    InMux I__5842 (
            .O(N__32024),
            .I(N__31981));
    InMux I__5841 (
            .O(N__32023),
            .I(N__31981));
    InMux I__5840 (
            .O(N__32022),
            .I(N__31970));
    InMux I__5839 (
            .O(N__32021),
            .I(N__31970));
    InMux I__5838 (
            .O(N__32020),
            .I(N__31970));
    InMux I__5837 (
            .O(N__32019),
            .I(N__31970));
    InMux I__5836 (
            .O(N__32018),
            .I(N__31970));
    InMux I__5835 (
            .O(N__32017),
            .I(N__31959));
    InMux I__5834 (
            .O(N__32016),
            .I(N__31959));
    InMux I__5833 (
            .O(N__32015),
            .I(N__31959));
    InMux I__5832 (
            .O(N__32014),
            .I(N__31959));
    InMux I__5831 (
            .O(N__32013),
            .I(N__31959));
    LocalMux I__5830 (
            .O(N__32010),
            .I(N__31956));
    InMux I__5829 (
            .O(N__32009),
            .I(N__31953));
    LocalMux I__5828 (
            .O(N__32006),
            .I(N__31950));
    InMux I__5827 (
            .O(N__32005),
            .I(N__31938));
    InMux I__5826 (
            .O(N__32004),
            .I(N__31938));
    InMux I__5825 (
            .O(N__32003),
            .I(N__31938));
    LocalMux I__5824 (
            .O(N__32000),
            .I(N__31935));
    LocalMux I__5823 (
            .O(N__31993),
            .I(N__31932));
    InMux I__5822 (
            .O(N__31992),
            .I(N__31929));
    LocalMux I__5821 (
            .O(N__31981),
            .I(N__31926));
    LocalMux I__5820 (
            .O(N__31970),
            .I(N__31923));
    LocalMux I__5819 (
            .O(N__31959),
            .I(N__31919));
    Span4Mux_v I__5818 (
            .O(N__31956),
            .I(N__31912));
    LocalMux I__5817 (
            .O(N__31953),
            .I(N__31912));
    Span4Mux_v I__5816 (
            .O(N__31950),
            .I(N__31912));
    InMux I__5815 (
            .O(N__31949),
            .I(N__31901));
    InMux I__5814 (
            .O(N__31948),
            .I(N__31901));
    InMux I__5813 (
            .O(N__31947),
            .I(N__31901));
    InMux I__5812 (
            .O(N__31946),
            .I(N__31901));
    InMux I__5811 (
            .O(N__31945),
            .I(N__31901));
    LocalMux I__5810 (
            .O(N__31938),
            .I(N__31894));
    Span4Mux_v I__5809 (
            .O(N__31935),
            .I(N__31894));
    Span4Mux_v I__5808 (
            .O(N__31932),
            .I(N__31894));
    LocalMux I__5807 (
            .O(N__31929),
            .I(N__31887));
    Span4Mux_v I__5806 (
            .O(N__31926),
            .I(N__31887));
    Span4Mux_h I__5805 (
            .O(N__31923),
            .I(N__31887));
    InMux I__5804 (
            .O(N__31922),
            .I(N__31884));
    Span4Mux_v I__5803 (
            .O(N__31919),
            .I(N__31879));
    Span4Mux_h I__5802 (
            .O(N__31912),
            .I(N__31879));
    LocalMux I__5801 (
            .O(N__31901),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__5800 (
            .O(N__31894),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__5799 (
            .O(N__31887),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__5798 (
            .O(N__31884),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__5797 (
            .O(N__31879),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    CascadeMux I__5796 (
            .O(N__31868),
            .I(N__31865));
    InMux I__5795 (
            .O(N__31865),
            .I(N__31861));
    CascadeMux I__5794 (
            .O(N__31864),
            .I(N__31858));
    LocalMux I__5793 (
            .O(N__31861),
            .I(N__31853));
    InMux I__5792 (
            .O(N__31858),
            .I(N__31850));
    InMux I__5791 (
            .O(N__31857),
            .I(N__31847));
    InMux I__5790 (
            .O(N__31856),
            .I(N__31844));
    Span4Mux_h I__5789 (
            .O(N__31853),
            .I(N__31838));
    LocalMux I__5788 (
            .O(N__31850),
            .I(N__31838));
    LocalMux I__5787 (
            .O(N__31847),
            .I(N__31833));
    LocalMux I__5786 (
            .O(N__31844),
            .I(N__31833));
    InMux I__5785 (
            .O(N__31843),
            .I(N__31830));
    Span4Mux_h I__5784 (
            .O(N__31838),
            .I(N__31827));
    Span12Mux_s11_h I__5783 (
            .O(N__31833),
            .I(N__31824));
    LocalMux I__5782 (
            .O(N__31830),
            .I(N__31821));
    Odrv4 I__5781 (
            .O(N__31827),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__5780 (
            .O(N__31824),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__5779 (
            .O(N__31821),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__5778 (
            .O(N__31814),
            .I(N__31811));
    LocalMux I__5777 (
            .O(N__31811),
            .I(N__31808));
    Span4Mux_h I__5776 (
            .O(N__31808),
            .I(N__31805));
    Span4Mux_h I__5775 (
            .O(N__31805),
            .I(N__31802));
    Odrv4 I__5774 (
            .O(N__31802),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__5773 (
            .O(N__31799),
            .I(N__31791));
    CascadeMux I__5772 (
            .O(N__31798),
            .I(N__31787));
    CascadeMux I__5771 (
            .O(N__31797),
            .I(N__31783));
    CascadeMux I__5770 (
            .O(N__31796),
            .I(N__31779));
    InMux I__5769 (
            .O(N__31795),
            .I(N__31761));
    InMux I__5768 (
            .O(N__31794),
            .I(N__31761));
    InMux I__5767 (
            .O(N__31791),
            .I(N__31761));
    InMux I__5766 (
            .O(N__31790),
            .I(N__31761));
    InMux I__5765 (
            .O(N__31787),
            .I(N__31761));
    InMux I__5764 (
            .O(N__31786),
            .I(N__31761));
    InMux I__5763 (
            .O(N__31783),
            .I(N__31761));
    InMux I__5762 (
            .O(N__31782),
            .I(N__31761));
    InMux I__5761 (
            .O(N__31779),
            .I(N__31752));
    InMux I__5760 (
            .O(N__31778),
            .I(N__31752));
    LocalMux I__5759 (
            .O(N__31761),
            .I(N__31749));
    CascadeMux I__5758 (
            .O(N__31760),
            .I(N__31746));
    CascadeMux I__5757 (
            .O(N__31759),
            .I(N__31742));
    CascadeMux I__5756 (
            .O(N__31758),
            .I(N__31738));
    CascadeMux I__5755 (
            .O(N__31757),
            .I(N__31734));
    LocalMux I__5754 (
            .O(N__31752),
            .I(N__31730));
    Span4Mux_v I__5753 (
            .O(N__31749),
            .I(N__31727));
    InMux I__5752 (
            .O(N__31746),
            .I(N__31710));
    InMux I__5751 (
            .O(N__31745),
            .I(N__31710));
    InMux I__5750 (
            .O(N__31742),
            .I(N__31710));
    InMux I__5749 (
            .O(N__31741),
            .I(N__31710));
    InMux I__5748 (
            .O(N__31738),
            .I(N__31710));
    InMux I__5747 (
            .O(N__31737),
            .I(N__31710));
    InMux I__5746 (
            .O(N__31734),
            .I(N__31710));
    InMux I__5745 (
            .O(N__31733),
            .I(N__31710));
    Span4Mux_h I__5744 (
            .O(N__31730),
            .I(N__31707));
    Span4Mux_h I__5743 (
            .O(N__31727),
            .I(N__31704));
    LocalMux I__5742 (
            .O(N__31710),
            .I(N__31701));
    Span4Mux_h I__5741 (
            .O(N__31707),
            .I(N__31698));
    Odrv4 I__5740 (
            .O(N__31704),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    Odrv12 I__5739 (
            .O(N__31701),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    Odrv4 I__5738 (
            .O(N__31698),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__5737 (
            .O(N__31691),
            .I(N__31688));
    LocalMux I__5736 (
            .O(N__31688),
            .I(N__31685));
    Span4Mux_v I__5735 (
            .O(N__31685),
            .I(N__31682));
    Span4Mux_v I__5734 (
            .O(N__31682),
            .I(N__31677));
    InMux I__5733 (
            .O(N__31681),
            .I(N__31672));
    InMux I__5732 (
            .O(N__31680),
            .I(N__31672));
    Sp12to4 I__5731 (
            .O(N__31677),
            .I(N__31667));
    LocalMux I__5730 (
            .O(N__31672),
            .I(N__31667));
    Span12Mux_h I__5729 (
            .O(N__31667),
            .I(N__31664));
    Span12Mux_v I__5728 (
            .O(N__31664),
            .I(N__31661));
    Odrv12 I__5727 (
            .O(N__31661),
            .I(il_max_comp2_c));
    InMux I__5726 (
            .O(N__31658),
            .I(N__31655));
    LocalMux I__5725 (
            .O(N__31655),
            .I(N__31651));
    InMux I__5724 (
            .O(N__31654),
            .I(N__31646));
    Span4Mux_h I__5723 (
            .O(N__31651),
            .I(N__31643));
    InMux I__5722 (
            .O(N__31650),
            .I(N__31640));
    InMux I__5721 (
            .O(N__31649),
            .I(N__31637));
    LocalMux I__5720 (
            .O(N__31646),
            .I(N__31634));
    Span4Mux_v I__5719 (
            .O(N__31643),
            .I(N__31631));
    LocalMux I__5718 (
            .O(N__31640),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__5717 (
            .O(N__31637),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__5716 (
            .O(N__31634),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__5715 (
            .O(N__31631),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    InMux I__5714 (
            .O(N__31622),
            .I(N__31619));
    LocalMux I__5713 (
            .O(N__31619),
            .I(N__31616));
    Odrv4 I__5712 (
            .O(N__31616),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt24 ));
    CascadeMux I__5711 (
            .O(N__31613),
            .I(N__31610));
    InMux I__5710 (
            .O(N__31610),
            .I(N__31607));
    LocalMux I__5709 (
            .O(N__31607),
            .I(N__31604));
    Odrv4 I__5708 (
            .O(N__31604),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ));
    InMux I__5707 (
            .O(N__31601),
            .I(N__31598));
    LocalMux I__5706 (
            .O(N__31598),
            .I(N__31595));
    Odrv4 I__5705 (
            .O(N__31595),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ));
    CascadeMux I__5704 (
            .O(N__31592),
            .I(N__31589));
    InMux I__5703 (
            .O(N__31589),
            .I(N__31586));
    LocalMux I__5702 (
            .O(N__31586),
            .I(N__31583));
    Span4Mux_h I__5701 (
            .O(N__31583),
            .I(N__31580));
    Span4Mux_h I__5700 (
            .O(N__31580),
            .I(N__31577));
    Odrv4 I__5699 (
            .O(N__31577),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt26 ));
    InMux I__5698 (
            .O(N__31574),
            .I(N__31571));
    LocalMux I__5697 (
            .O(N__31571),
            .I(N__31568));
    Span4Mux_h I__5696 (
            .O(N__31568),
            .I(N__31565));
    Odrv4 I__5695 (
            .O(N__31565),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ));
    CascadeMux I__5694 (
            .O(N__31562),
            .I(N__31559));
    InMux I__5693 (
            .O(N__31559),
            .I(N__31556));
    LocalMux I__5692 (
            .O(N__31556),
            .I(N__31553));
    Span4Mux_h I__5691 (
            .O(N__31553),
            .I(N__31550));
    Odrv4 I__5690 (
            .O(N__31550),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt28 ));
    InMux I__5689 (
            .O(N__31547),
            .I(N__31544));
    LocalMux I__5688 (
            .O(N__31544),
            .I(N__31541));
    Span4Mux_v I__5687 (
            .O(N__31541),
            .I(N__31538));
    Odrv4 I__5686 (
            .O(N__31538),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ));
    CascadeMux I__5685 (
            .O(N__31535),
            .I(N__31532));
    InMux I__5684 (
            .O(N__31532),
            .I(N__31528));
    CascadeMux I__5683 (
            .O(N__31531),
            .I(N__31525));
    LocalMux I__5682 (
            .O(N__31528),
            .I(N__31522));
    InMux I__5681 (
            .O(N__31525),
            .I(N__31519));
    Span4Mux_v I__5680 (
            .O(N__31522),
            .I(N__31514));
    LocalMux I__5679 (
            .O(N__31519),
            .I(N__31514));
    Odrv4 I__5678 (
            .O(N__31514),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    InMux I__5677 (
            .O(N__31511),
            .I(N__31508));
    LocalMux I__5676 (
            .O(N__31508),
            .I(N__31505));
    Sp12to4 I__5675 (
            .O(N__31505),
            .I(N__31502));
    Odrv12 I__5674 (
            .O(N__31502),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ));
    InMux I__5673 (
            .O(N__31499),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ));
    InMux I__5672 (
            .O(N__31496),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    InMux I__5671 (
            .O(N__31493),
            .I(N__31490));
    LocalMux I__5670 (
            .O(N__31490),
            .I(N__31486));
    InMux I__5669 (
            .O(N__31489),
            .I(N__31482));
    Span4Mux_h I__5668 (
            .O(N__31486),
            .I(N__31479));
    InMux I__5667 (
            .O(N__31485),
            .I(N__31476));
    LocalMux I__5666 (
            .O(N__31482),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    Odrv4 I__5665 (
            .O(N__31479),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    LocalMux I__5664 (
            .O(N__31476),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    CascadeMux I__5663 (
            .O(N__31469),
            .I(N__31466));
    InMux I__5662 (
            .O(N__31466),
            .I(N__31462));
    InMux I__5661 (
            .O(N__31465),
            .I(N__31458));
    LocalMux I__5660 (
            .O(N__31462),
            .I(N__31455));
    InMux I__5659 (
            .O(N__31461),
            .I(N__31452));
    LocalMux I__5658 (
            .O(N__31458),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    Odrv4 I__5657 (
            .O(N__31455),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    LocalMux I__5656 (
            .O(N__31452),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    InMux I__5655 (
            .O(N__31445),
            .I(N__31442));
    LocalMux I__5654 (
            .O(N__31442),
            .I(N__31437));
    CascadeMux I__5653 (
            .O(N__31441),
            .I(N__31434));
    InMux I__5652 (
            .O(N__31440),
            .I(N__31431));
    Span4Mux_v I__5651 (
            .O(N__31437),
            .I(N__31428));
    InMux I__5650 (
            .O(N__31434),
            .I(N__31425));
    LocalMux I__5649 (
            .O(N__31431),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    Odrv4 I__5648 (
            .O(N__31428),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    LocalMux I__5647 (
            .O(N__31425),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    InMux I__5646 (
            .O(N__31418),
            .I(N__31415));
    LocalMux I__5645 (
            .O(N__31415),
            .I(N__31411));
    InMux I__5644 (
            .O(N__31414),
            .I(N__31407));
    Span4Mux_h I__5643 (
            .O(N__31411),
            .I(N__31404));
    InMux I__5642 (
            .O(N__31410),
            .I(N__31401));
    LocalMux I__5641 (
            .O(N__31407),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    Odrv4 I__5640 (
            .O(N__31404),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    LocalMux I__5639 (
            .O(N__31401),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    CascadeMux I__5638 (
            .O(N__31394),
            .I(N__31391));
    InMux I__5637 (
            .O(N__31391),
            .I(N__31388));
    LocalMux I__5636 (
            .O(N__31388),
            .I(N__31385));
    Span4Mux_v I__5635 (
            .O(N__31385),
            .I(N__31382));
    Odrv4 I__5634 (
            .O(N__31382),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    InMux I__5633 (
            .O(N__31379),
            .I(N__31375));
    InMux I__5632 (
            .O(N__31378),
            .I(N__31372));
    LocalMux I__5631 (
            .O(N__31375),
            .I(N__31369));
    LocalMux I__5630 (
            .O(N__31372),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv12 I__5629 (
            .O(N__31369),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__5628 (
            .O(N__31364),
            .I(N__31361));
    LocalMux I__5627 (
            .O(N__31361),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__5626 (
            .O(N__31358),
            .I(N__31354));
    InMux I__5625 (
            .O(N__31357),
            .I(N__31351));
    LocalMux I__5624 (
            .O(N__31354),
            .I(N__31348));
    LocalMux I__5623 (
            .O(N__31351),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv12 I__5622 (
            .O(N__31348),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__5621 (
            .O(N__31343),
            .I(N__31340));
    LocalMux I__5620 (
            .O(N__31340),
            .I(N__31337));
    Span4Mux_v I__5619 (
            .O(N__31337),
            .I(N__31334));
    Odrv4 I__5618 (
            .O(N__31334),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__5617 (
            .O(N__31331),
            .I(N__31328));
    InMux I__5616 (
            .O(N__31328),
            .I(N__31325));
    LocalMux I__5615 (
            .O(N__31325),
            .I(N__31322));
    Odrv4 I__5614 (
            .O(N__31322),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__5613 (
            .O(N__31319),
            .I(N__31315));
    InMux I__5612 (
            .O(N__31318),
            .I(N__31312));
    LocalMux I__5611 (
            .O(N__31315),
            .I(N__31309));
    LocalMux I__5610 (
            .O(N__31312),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv12 I__5609 (
            .O(N__31309),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__5608 (
            .O(N__31304),
            .I(N__31301));
    InMux I__5607 (
            .O(N__31301),
            .I(N__31298));
    LocalMux I__5606 (
            .O(N__31298),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__5605 (
            .O(N__31295),
            .I(N__31291));
    InMux I__5604 (
            .O(N__31294),
            .I(N__31288));
    LocalMux I__5603 (
            .O(N__31291),
            .I(N__31285));
    LocalMux I__5602 (
            .O(N__31288),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv12 I__5601 (
            .O(N__31285),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__5600 (
            .O(N__31280),
            .I(N__31277));
    LocalMux I__5599 (
            .O(N__31277),
            .I(N__31274));
    Odrv4 I__5598 (
            .O(N__31274),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__5597 (
            .O(N__31271),
            .I(N__31268));
    InMux I__5596 (
            .O(N__31268),
            .I(N__31265));
    LocalMux I__5595 (
            .O(N__31265),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__5594 (
            .O(N__31262),
            .I(N__31259));
    LocalMux I__5593 (
            .O(N__31259),
            .I(N__31256));
    Span4Mux_v I__5592 (
            .O(N__31256),
            .I(N__31253));
    Odrv4 I__5591 (
            .O(N__31253),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    CascadeMux I__5590 (
            .O(N__31250),
            .I(N__31247));
    InMux I__5589 (
            .O(N__31247),
            .I(N__31244));
    LocalMux I__5588 (
            .O(N__31244),
            .I(N__31241));
    Span4Mux_h I__5587 (
            .O(N__31241),
            .I(N__31238));
    Span4Mux_v I__5586 (
            .O(N__31238),
            .I(N__31235));
    Odrv4 I__5585 (
            .O(N__31235),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__5584 (
            .O(N__31232),
            .I(N__31229));
    LocalMux I__5583 (
            .O(N__31229),
            .I(N__31226));
    Odrv4 I__5582 (
            .O(N__31226),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ));
    CascadeMux I__5581 (
            .O(N__31223),
            .I(N__31220));
    InMux I__5580 (
            .O(N__31220),
            .I(N__31217));
    LocalMux I__5579 (
            .O(N__31217),
            .I(N__31214));
    Span4Mux_v I__5578 (
            .O(N__31214),
            .I(N__31211));
    Odrv4 I__5577 (
            .O(N__31211),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt20 ));
    InMux I__5576 (
            .O(N__31208),
            .I(N__31205));
    LocalMux I__5575 (
            .O(N__31205),
            .I(N__31202));
    Odrv12 I__5574 (
            .O(N__31202),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ));
    CascadeMux I__5573 (
            .O(N__31199),
            .I(N__31196));
    InMux I__5572 (
            .O(N__31196),
            .I(N__31193));
    LocalMux I__5571 (
            .O(N__31193),
            .I(N__31190));
    Odrv12 I__5570 (
            .O(N__31190),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt22 ));
    InMux I__5569 (
            .O(N__31187),
            .I(N__31183));
    InMux I__5568 (
            .O(N__31186),
            .I(N__31180));
    LocalMux I__5567 (
            .O(N__31183),
            .I(N__31177));
    LocalMux I__5566 (
            .O(N__31180),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv12 I__5565 (
            .O(N__31177),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__5564 (
            .O(N__31172),
            .I(N__31169));
    LocalMux I__5563 (
            .O(N__31169),
            .I(N__31166));
    Span4Mux_v I__5562 (
            .O(N__31166),
            .I(N__31163));
    Span4Mux_v I__5561 (
            .O(N__31163),
            .I(N__31160));
    Odrv4 I__5560 (
            .O(N__31160),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__5559 (
            .O(N__31157),
            .I(N__31154));
    InMux I__5558 (
            .O(N__31154),
            .I(N__31151));
    LocalMux I__5557 (
            .O(N__31151),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__5556 (
            .O(N__31148),
            .I(N__31144));
    InMux I__5555 (
            .O(N__31147),
            .I(N__31141));
    LocalMux I__5554 (
            .O(N__31144),
            .I(N__31138));
    LocalMux I__5553 (
            .O(N__31141),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv12 I__5552 (
            .O(N__31138),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__5551 (
            .O(N__31133),
            .I(N__31130));
    LocalMux I__5550 (
            .O(N__31130),
            .I(N__31127));
    Span4Mux_v I__5549 (
            .O(N__31127),
            .I(N__31124));
    Odrv4 I__5548 (
            .O(N__31124),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__5547 (
            .O(N__31121),
            .I(N__31118));
    InMux I__5546 (
            .O(N__31118),
            .I(N__31115));
    LocalMux I__5545 (
            .O(N__31115),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__5544 (
            .O(N__31112),
            .I(N__31109));
    LocalMux I__5543 (
            .O(N__31109),
            .I(N__31106));
    Span4Mux_v I__5542 (
            .O(N__31106),
            .I(N__31103));
    Odrv4 I__5541 (
            .O(N__31103),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__5540 (
            .O(N__31100),
            .I(N__31097));
    LocalMux I__5539 (
            .O(N__31097),
            .I(N__31093));
    InMux I__5538 (
            .O(N__31096),
            .I(N__31090));
    Span4Mux_v I__5537 (
            .O(N__31093),
            .I(N__31087));
    LocalMux I__5536 (
            .O(N__31090),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__5535 (
            .O(N__31087),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__5534 (
            .O(N__31082),
            .I(N__31079));
    InMux I__5533 (
            .O(N__31079),
            .I(N__31076));
    LocalMux I__5532 (
            .O(N__31076),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__5531 (
            .O(N__31073),
            .I(N__31070));
    LocalMux I__5530 (
            .O(N__31070),
            .I(N__31067));
    Span4Mux_v I__5529 (
            .O(N__31067),
            .I(N__31064));
    Odrv4 I__5528 (
            .O(N__31064),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    InMux I__5527 (
            .O(N__31061),
            .I(N__31058));
    LocalMux I__5526 (
            .O(N__31058),
            .I(N__31054));
    InMux I__5525 (
            .O(N__31057),
            .I(N__31051));
    Span4Mux_v I__5524 (
            .O(N__31054),
            .I(N__31048));
    LocalMux I__5523 (
            .O(N__31051),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__5522 (
            .O(N__31048),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__5521 (
            .O(N__31043),
            .I(N__31040));
    InMux I__5520 (
            .O(N__31040),
            .I(N__31037));
    LocalMux I__5519 (
            .O(N__31037),
            .I(N__31034));
    Odrv12 I__5518 (
            .O(N__31034),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__5517 (
            .O(N__31031),
            .I(N__31028));
    LocalMux I__5516 (
            .O(N__31028),
            .I(N__31025));
    Span4Mux_v I__5515 (
            .O(N__31025),
            .I(N__31022));
    Odrv4 I__5514 (
            .O(N__31022),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__5513 (
            .O(N__31019),
            .I(N__31015));
    InMux I__5512 (
            .O(N__31018),
            .I(N__31012));
    LocalMux I__5511 (
            .O(N__31015),
            .I(N__31009));
    LocalMux I__5510 (
            .O(N__31012),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv12 I__5509 (
            .O(N__31009),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__5508 (
            .O(N__31004),
            .I(N__31001));
    InMux I__5507 (
            .O(N__31001),
            .I(N__30998));
    LocalMux I__5506 (
            .O(N__30998),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__5505 (
            .O(N__30995),
            .I(N__30991));
    InMux I__5504 (
            .O(N__30994),
            .I(N__30988));
    LocalMux I__5503 (
            .O(N__30991),
            .I(N__30985));
    LocalMux I__5502 (
            .O(N__30988),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv12 I__5501 (
            .O(N__30985),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__5500 (
            .O(N__30980),
            .I(N__30977));
    InMux I__5499 (
            .O(N__30977),
            .I(N__30974));
    LocalMux I__5498 (
            .O(N__30974),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__5497 (
            .O(N__30971),
            .I(N__30968));
    LocalMux I__5496 (
            .O(N__30968),
            .I(N__30965));
    Span4Mux_h I__5495 (
            .O(N__30965),
            .I(N__30962));
    Span4Mux_v I__5494 (
            .O(N__30962),
            .I(N__30959));
    Odrv4 I__5493 (
            .O(N__30959),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__5492 (
            .O(N__30956),
            .I(N__30952));
    InMux I__5491 (
            .O(N__30955),
            .I(N__30949));
    LocalMux I__5490 (
            .O(N__30952),
            .I(N__30946));
    LocalMux I__5489 (
            .O(N__30949),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv12 I__5488 (
            .O(N__30946),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    CascadeMux I__5487 (
            .O(N__30941),
            .I(N__30938));
    InMux I__5486 (
            .O(N__30938),
            .I(N__30935));
    LocalMux I__5485 (
            .O(N__30935),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__5484 (
            .O(N__30932),
            .I(N__30925));
    InMux I__5483 (
            .O(N__30931),
            .I(N__30925));
    InMux I__5482 (
            .O(N__30930),
            .I(N__30922));
    LocalMux I__5481 (
            .O(N__30925),
            .I(N__30919));
    LocalMux I__5480 (
            .O(N__30922),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__5479 (
            .O(N__30919),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__5478 (
            .O(N__30914),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    CascadeMux I__5477 (
            .O(N__30911),
            .I(N__30908));
    InMux I__5476 (
            .O(N__30908),
            .I(N__30898));
    InMux I__5475 (
            .O(N__30907),
            .I(N__30898));
    InMux I__5474 (
            .O(N__30906),
            .I(N__30898));
    InMux I__5473 (
            .O(N__30905),
            .I(N__30895));
    LocalMux I__5472 (
            .O(N__30898),
            .I(N__30892));
    LocalMux I__5471 (
            .O(N__30895),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__5470 (
            .O(N__30892),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__5469 (
            .O(N__30887),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__5468 (
            .O(N__30884),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__5467 (
            .O(N__30881),
            .I(N__30871));
    InMux I__5466 (
            .O(N__30880),
            .I(N__30871));
    InMux I__5465 (
            .O(N__30879),
            .I(N__30871));
    InMux I__5464 (
            .O(N__30878),
            .I(N__30868));
    LocalMux I__5463 (
            .O(N__30871),
            .I(N__30865));
    LocalMux I__5462 (
            .O(N__30868),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__5461 (
            .O(N__30865),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__5460 (
            .O(N__30860),
            .I(N__30857));
    LocalMux I__5459 (
            .O(N__30857),
            .I(N__30853));
    InMux I__5458 (
            .O(N__30856),
            .I(N__30850));
    Odrv12 I__5457 (
            .O(N__30853),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__5456 (
            .O(N__30850),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    InMux I__5455 (
            .O(N__30845),
            .I(N__30842));
    LocalMux I__5454 (
            .O(N__30842),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__5453 (
            .O(N__30839),
            .I(N__30836));
    InMux I__5452 (
            .O(N__30836),
            .I(N__30832));
    CascadeMux I__5451 (
            .O(N__30835),
            .I(N__30829));
    LocalMux I__5450 (
            .O(N__30832),
            .I(N__30826));
    InMux I__5449 (
            .O(N__30829),
            .I(N__30822));
    Span4Mux_h I__5448 (
            .O(N__30826),
            .I(N__30819));
    InMux I__5447 (
            .O(N__30825),
            .I(N__30816));
    LocalMux I__5446 (
            .O(N__30822),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__5445 (
            .O(N__30819),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__5444 (
            .O(N__30816),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__5443 (
            .O(N__30809),
            .I(N__30806));
    InMux I__5442 (
            .O(N__30806),
            .I(N__30803));
    LocalMux I__5441 (
            .O(N__30803),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__5440 (
            .O(N__30800),
            .I(N__30797));
    LocalMux I__5439 (
            .O(N__30797),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__5438 (
            .O(N__30794),
            .I(N__30790));
    InMux I__5437 (
            .O(N__30793),
            .I(N__30787));
    LocalMux I__5436 (
            .O(N__30790),
            .I(N__30784));
    LocalMux I__5435 (
            .O(N__30787),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv12 I__5434 (
            .O(N__30784),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    CascadeMux I__5433 (
            .O(N__30779),
            .I(N__30776));
    InMux I__5432 (
            .O(N__30776),
            .I(N__30773));
    LocalMux I__5431 (
            .O(N__30773),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__5430 (
            .O(N__30770),
            .I(N__30767));
    LocalMux I__5429 (
            .O(N__30767),
            .I(N__30763));
    InMux I__5428 (
            .O(N__30766),
            .I(N__30760));
    Span4Mux_v I__5427 (
            .O(N__30763),
            .I(N__30757));
    LocalMux I__5426 (
            .O(N__30760),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__5425 (
            .O(N__30757),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__5424 (
            .O(N__30752),
            .I(N__30749));
    LocalMux I__5423 (
            .O(N__30749),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__5422 (
            .O(N__30746),
            .I(N__30743));
    InMux I__5421 (
            .O(N__30743),
            .I(N__30740));
    LocalMux I__5420 (
            .O(N__30740),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__5419 (
            .O(N__30737),
            .I(N__30734));
    InMux I__5418 (
            .O(N__30734),
            .I(N__30731));
    LocalMux I__5417 (
            .O(N__30731),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__5416 (
            .O(N__30728),
            .I(N__30724));
    InMux I__5415 (
            .O(N__30727),
            .I(N__30721));
    LocalMux I__5414 (
            .O(N__30724),
            .I(N__30718));
    LocalMux I__5413 (
            .O(N__30721),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv12 I__5412 (
            .O(N__30718),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__5411 (
            .O(N__30713),
            .I(N__30710));
    LocalMux I__5410 (
            .O(N__30710),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__5409 (
            .O(N__30707),
            .I(N__30703));
    InMux I__5408 (
            .O(N__30706),
            .I(N__30699));
    InMux I__5407 (
            .O(N__30703),
            .I(N__30694));
    InMux I__5406 (
            .O(N__30702),
            .I(N__30694));
    LocalMux I__5405 (
            .O(N__30699),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    LocalMux I__5404 (
            .O(N__30694),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__5403 (
            .O(N__30689),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__5402 (
            .O(N__30686),
            .I(N__30683));
    InMux I__5401 (
            .O(N__30683),
            .I(N__30677));
    InMux I__5400 (
            .O(N__30682),
            .I(N__30677));
    LocalMux I__5399 (
            .O(N__30677),
            .I(N__30673));
    InMux I__5398 (
            .O(N__30676),
            .I(N__30670));
    Span4Mux_h I__5397 (
            .O(N__30673),
            .I(N__30667));
    LocalMux I__5396 (
            .O(N__30670),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__5395 (
            .O(N__30667),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__5394 (
            .O(N__30662),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__5393 (
            .O(N__30659),
            .I(N__30652));
    InMux I__5392 (
            .O(N__30658),
            .I(N__30652));
    InMux I__5391 (
            .O(N__30657),
            .I(N__30649));
    LocalMux I__5390 (
            .O(N__30652),
            .I(N__30646));
    LocalMux I__5389 (
            .O(N__30649),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv12 I__5388 (
            .O(N__30646),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__5387 (
            .O(N__30641),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__5386 (
            .O(N__30638),
            .I(N__30631));
    InMux I__5385 (
            .O(N__30637),
            .I(N__30631));
    InMux I__5384 (
            .O(N__30636),
            .I(N__30628));
    LocalMux I__5383 (
            .O(N__30631),
            .I(N__30625));
    LocalMux I__5382 (
            .O(N__30628),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__5381 (
            .O(N__30625),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__5380 (
            .O(N__30620),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__5379 (
            .O(N__30617),
            .I(N__30612));
    InMux I__5378 (
            .O(N__30616),
            .I(N__30609));
    InMux I__5377 (
            .O(N__30615),
            .I(N__30606));
    LocalMux I__5376 (
            .O(N__30612),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    LocalMux I__5375 (
            .O(N__30609),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    LocalMux I__5374 (
            .O(N__30606),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__5373 (
            .O(N__30599),
            .I(bfn_11_12_0_));
    CascadeMux I__5372 (
            .O(N__30596),
            .I(N__30593));
    InMux I__5371 (
            .O(N__30593),
            .I(N__30589));
    CascadeMux I__5370 (
            .O(N__30592),
            .I(N__30585));
    LocalMux I__5369 (
            .O(N__30589),
            .I(N__30582));
    InMux I__5368 (
            .O(N__30588),
            .I(N__30579));
    InMux I__5367 (
            .O(N__30585),
            .I(N__30576));
    Span4Mux_h I__5366 (
            .O(N__30582),
            .I(N__30573));
    LocalMux I__5365 (
            .O(N__30579),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__5364 (
            .O(N__30576),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv4 I__5363 (
            .O(N__30573),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__5362 (
            .O(N__30566),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__5361 (
            .O(N__30563),
            .I(N__30559));
    InMux I__5360 (
            .O(N__30562),
            .I(N__30555));
    LocalMux I__5359 (
            .O(N__30559),
            .I(N__30552));
    InMux I__5358 (
            .O(N__30558),
            .I(N__30549));
    LocalMux I__5357 (
            .O(N__30555),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__5356 (
            .O(N__30552),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__5355 (
            .O(N__30549),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__5354 (
            .O(N__30542),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    CascadeMux I__5353 (
            .O(N__30539),
            .I(N__30535));
    InMux I__5352 (
            .O(N__30538),
            .I(N__30529));
    InMux I__5351 (
            .O(N__30535),
            .I(N__30529));
    InMux I__5350 (
            .O(N__30534),
            .I(N__30526));
    LocalMux I__5349 (
            .O(N__30529),
            .I(N__30523));
    LocalMux I__5348 (
            .O(N__30526),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__5347 (
            .O(N__30523),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__5346 (
            .O(N__30518),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__5345 (
            .O(N__30515),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__5344 (
            .O(N__30512),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__5343 (
            .O(N__30509),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__5342 (
            .O(N__30506),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__5341 (
            .O(N__30503),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__5340 (
            .O(N__30500),
            .I(bfn_11_11_0_));
    CascadeMux I__5339 (
            .O(N__30497),
            .I(N__30493));
    InMux I__5338 (
            .O(N__30496),
            .I(N__30489));
    InMux I__5337 (
            .O(N__30493),
            .I(N__30484));
    InMux I__5336 (
            .O(N__30492),
            .I(N__30484));
    LocalMux I__5335 (
            .O(N__30489),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__5334 (
            .O(N__30484),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__5333 (
            .O(N__30479),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__5332 (
            .O(N__30476),
            .I(N__30471));
    InMux I__5331 (
            .O(N__30475),
            .I(N__30466));
    InMux I__5330 (
            .O(N__30474),
            .I(N__30466));
    LocalMux I__5329 (
            .O(N__30471),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__5328 (
            .O(N__30466),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__5327 (
            .O(N__30461),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__5326 (
            .O(N__30458),
            .I(N__30453));
    InMux I__5325 (
            .O(N__30457),
            .I(N__30448));
    InMux I__5324 (
            .O(N__30456),
            .I(N__30448));
    LocalMux I__5323 (
            .O(N__30453),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    LocalMux I__5322 (
            .O(N__30448),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__5321 (
            .O(N__30443),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    CascadeMux I__5320 (
            .O(N__30440),
            .I(N__30437));
    InMux I__5319 (
            .O(N__30437),
            .I(N__30434));
    LocalMux I__5318 (
            .O(N__30434),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ));
    InMux I__5317 (
            .O(N__30431),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__5316 (
            .O(N__30428),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__5315 (
            .O(N__30425),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__5314 (
            .O(N__30422),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__5313 (
            .O(N__30419),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__5312 (
            .O(N__30416),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__5311 (
            .O(N__30413),
            .I(bfn_11_10_0_));
    InMux I__5310 (
            .O(N__30410),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__5309 (
            .O(N__30407),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__5308 (
            .O(N__30404),
            .I(N__30400));
    InMux I__5307 (
            .O(N__30403),
            .I(N__30396));
    LocalMux I__5306 (
            .O(N__30400),
            .I(N__30393));
    InMux I__5305 (
            .O(N__30399),
            .I(N__30390));
    LocalMux I__5304 (
            .O(N__30396),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    Odrv12 I__5303 (
            .O(N__30393),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    LocalMux I__5302 (
            .O(N__30390),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__5301 (
            .O(N__30383),
            .I(N__30379));
    InMux I__5300 (
            .O(N__30382),
            .I(N__30376));
    LocalMux I__5299 (
            .O(N__30379),
            .I(N__30372));
    LocalMux I__5298 (
            .O(N__30376),
            .I(N__30369));
    InMux I__5297 (
            .O(N__30375),
            .I(N__30365));
    Span4Mux_h I__5296 (
            .O(N__30372),
            .I(N__30360));
    Span4Mux_h I__5295 (
            .O(N__30369),
            .I(N__30360));
    InMux I__5294 (
            .O(N__30368),
            .I(N__30357));
    LocalMux I__5293 (
            .O(N__30365),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv4 I__5292 (
            .O(N__30360),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__5291 (
            .O(N__30357),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__5290 (
            .O(N__30350),
            .I(N__30347));
    LocalMux I__5289 (
            .O(N__30347),
            .I(N__30344));
    Odrv4 I__5288 (
            .O(N__30344),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df30 ));
    CascadeMux I__5287 (
            .O(N__30341),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__5286 (
            .O(N__30338),
            .I(N__30332));
    InMux I__5285 (
            .O(N__30337),
            .I(N__30332));
    LocalMux I__5284 (
            .O(N__30332),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    CascadeMux I__5283 (
            .O(N__30329),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ));
    InMux I__5282 (
            .O(N__30326),
            .I(N__30323));
    LocalMux I__5281 (
            .O(N__30323),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    InMux I__5280 (
            .O(N__30320),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__5279 (
            .O(N__30317),
            .I(N__30313));
    CascadeMux I__5278 (
            .O(N__30316),
            .I(N__30309));
    InMux I__5277 (
            .O(N__30313),
            .I(N__30302));
    InMux I__5276 (
            .O(N__30312),
            .I(N__30302));
    InMux I__5275 (
            .O(N__30309),
            .I(N__30302));
    LocalMux I__5274 (
            .O(N__30302),
            .I(N__30299));
    Odrv4 I__5273 (
            .O(N__30299),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ));
    InMux I__5272 (
            .O(N__30296),
            .I(N__30293));
    LocalMux I__5271 (
            .O(N__30293),
            .I(N__30290));
    Span4Mux_h I__5270 (
            .O(N__30290),
            .I(N__30287));
    Odrv4 I__5269 (
            .O(N__30287),
            .I(il_min_comp1_c));
    InMux I__5268 (
            .O(N__30284),
            .I(N__30281));
    LocalMux I__5267 (
            .O(N__30281),
            .I(il_max_comp1_D1));
    InMux I__5266 (
            .O(N__30278),
            .I(N__30275));
    LocalMux I__5265 (
            .O(N__30275),
            .I(N__30270));
    InMux I__5264 (
            .O(N__30274),
            .I(N__30267));
    InMux I__5263 (
            .O(N__30273),
            .I(N__30264));
    Span4Mux_h I__5262 (
            .O(N__30270),
            .I(N__30260));
    LocalMux I__5261 (
            .O(N__30267),
            .I(N__30257));
    LocalMux I__5260 (
            .O(N__30264),
            .I(N__30254));
    InMux I__5259 (
            .O(N__30263),
            .I(N__30251));
    Odrv4 I__5258 (
            .O(N__30260),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv4 I__5257 (
            .O(N__30257),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv4 I__5256 (
            .O(N__30254),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__5255 (
            .O(N__30251),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__5254 (
            .O(N__30242),
            .I(N__30239));
    LocalMux I__5253 (
            .O(N__30239),
            .I(N__30235));
    InMux I__5252 (
            .O(N__30238),
            .I(N__30231));
    Span4Mux_h I__5251 (
            .O(N__30235),
            .I(N__30228));
    InMux I__5250 (
            .O(N__30234),
            .I(N__30225));
    LocalMux I__5249 (
            .O(N__30231),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv4 I__5248 (
            .O(N__30228),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    LocalMux I__5247 (
            .O(N__30225),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    InMux I__5246 (
            .O(N__30218),
            .I(N__30215));
    LocalMux I__5245 (
            .O(N__30215),
            .I(N__30212));
    Span4Mux_v I__5244 (
            .O(N__30212),
            .I(N__30208));
    InMux I__5243 (
            .O(N__30211),
            .I(N__30205));
    Odrv4 I__5242 (
            .O(N__30208),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__5241 (
            .O(N__30205),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    CascadeMux I__5240 (
            .O(N__30200),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23_cascade_));
    CascadeMux I__5239 (
            .O(N__30197),
            .I(N__30192));
    InMux I__5238 (
            .O(N__30196),
            .I(N__30187));
    InMux I__5237 (
            .O(N__30195),
            .I(N__30187));
    InMux I__5236 (
            .O(N__30192),
            .I(N__30184));
    LocalMux I__5235 (
            .O(N__30187),
            .I(N__30181));
    LocalMux I__5234 (
            .O(N__30184),
            .I(N__30177));
    Span4Mux_v I__5233 (
            .O(N__30181),
            .I(N__30174));
    InMux I__5232 (
            .O(N__30180),
            .I(N__30171));
    Odrv4 I__5231 (
            .O(N__30177),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    Odrv4 I__5230 (
            .O(N__30174),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__5229 (
            .O(N__30171),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    CascadeMux I__5228 (
            .O(N__30164),
            .I(N__30161));
    InMux I__5227 (
            .O(N__30161),
            .I(N__30155));
    InMux I__5226 (
            .O(N__30160),
            .I(N__30155));
    LocalMux I__5225 (
            .O(N__30155),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    InMux I__5224 (
            .O(N__30152),
            .I(N__30148));
    InMux I__5223 (
            .O(N__30151),
            .I(N__30144));
    LocalMux I__5222 (
            .O(N__30148),
            .I(N__30141));
    InMux I__5221 (
            .O(N__30147),
            .I(N__30138));
    LocalMux I__5220 (
            .O(N__30144),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv12 I__5219 (
            .O(N__30141),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    LocalMux I__5218 (
            .O(N__30138),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    InMux I__5217 (
            .O(N__30131),
            .I(N__30127));
    InMux I__5216 (
            .O(N__30130),
            .I(N__30123));
    LocalMux I__5215 (
            .O(N__30127),
            .I(N__30120));
    InMux I__5214 (
            .O(N__30126),
            .I(N__30117));
    LocalMux I__5213 (
            .O(N__30123),
            .I(N__30114));
    Span4Mux_v I__5212 (
            .O(N__30120),
            .I(N__30108));
    LocalMux I__5211 (
            .O(N__30117),
            .I(N__30108));
    Span4Mux_h I__5210 (
            .O(N__30114),
            .I(N__30105));
    InMux I__5209 (
            .O(N__30113),
            .I(N__30102));
    Odrv4 I__5208 (
            .O(N__30108),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv4 I__5207 (
            .O(N__30105),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    LocalMux I__5206 (
            .O(N__30102),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__5205 (
            .O(N__30095),
            .I(N__30091));
    InMux I__5204 (
            .O(N__30094),
            .I(N__30086));
    LocalMux I__5203 (
            .O(N__30091),
            .I(N__30083));
    InMux I__5202 (
            .O(N__30090),
            .I(N__30080));
    InMux I__5201 (
            .O(N__30089),
            .I(N__30077));
    LocalMux I__5200 (
            .O(N__30086),
            .I(N__30073));
    Span4Mux_h I__5199 (
            .O(N__30083),
            .I(N__30070));
    LocalMux I__5198 (
            .O(N__30080),
            .I(N__30065));
    LocalMux I__5197 (
            .O(N__30077),
            .I(N__30065));
    InMux I__5196 (
            .O(N__30076),
            .I(N__30062));
    Span4Mux_v I__5195 (
            .O(N__30073),
            .I(N__30059));
    Span4Mux_v I__5194 (
            .O(N__30070),
            .I(N__30054));
    Span4Mux_h I__5193 (
            .O(N__30065),
            .I(N__30054));
    LocalMux I__5192 (
            .O(N__30062),
            .I(N__30051));
    Odrv4 I__5191 (
            .O(N__30059),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__5190 (
            .O(N__30054),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__5189 (
            .O(N__30051),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__5188 (
            .O(N__30044),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_31 ));
    CascadeMux I__5187 (
            .O(N__30041),
            .I(N__30038));
    InMux I__5186 (
            .O(N__30038),
            .I(N__30035));
    LocalMux I__5185 (
            .O(N__30035),
            .I(N__30032));
    Span4Mux_h I__5184 (
            .O(N__30032),
            .I(N__30029));
    Odrv4 I__5183 (
            .O(N__30029),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0 ));
    InMux I__5182 (
            .O(N__30026),
            .I(N__30021));
    InMux I__5181 (
            .O(N__30025),
            .I(N__30018));
    InMux I__5180 (
            .O(N__30024),
            .I(N__30015));
    LocalMux I__5179 (
            .O(N__30021),
            .I(N__30012));
    LocalMux I__5178 (
            .O(N__30018),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    LocalMux I__5177 (
            .O(N__30015),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    Odrv4 I__5176 (
            .O(N__30012),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    CascadeMux I__5175 (
            .O(N__30005),
            .I(N__30001));
    InMux I__5174 (
            .O(N__30004),
            .I(N__29997));
    InMux I__5173 (
            .O(N__30001),
            .I(N__29994));
    InMux I__5172 (
            .O(N__30000),
            .I(N__29991));
    LocalMux I__5171 (
            .O(N__29997),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    LocalMux I__5170 (
            .O(N__29994),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    LocalMux I__5169 (
            .O(N__29991),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    CascadeMux I__5168 (
            .O(N__29984),
            .I(N__29981));
    InMux I__5167 (
            .O(N__29981),
            .I(N__29978));
    LocalMux I__5166 (
            .O(N__29978),
            .I(N__29973));
    InMux I__5165 (
            .O(N__29977),
            .I(N__29970));
    InMux I__5164 (
            .O(N__29976),
            .I(N__29967));
    Span4Mux_h I__5163 (
            .O(N__29973),
            .I(N__29962));
    LocalMux I__5162 (
            .O(N__29970),
            .I(N__29957));
    LocalMux I__5161 (
            .O(N__29967),
            .I(N__29957));
    InMux I__5160 (
            .O(N__29966),
            .I(N__29952));
    InMux I__5159 (
            .O(N__29965),
            .I(N__29952));
    Odrv4 I__5158 (
            .O(N__29962),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv12 I__5157 (
            .O(N__29957),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__5156 (
            .O(N__29952),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__5155 (
            .O(N__29945),
            .I(N__29942));
    LocalMux I__5154 (
            .O(N__29942),
            .I(N__29939));
    Odrv4 I__5153 (
            .O(N__29939),
            .I(\current_shift_inst.PI_CTRL.integrator_i_22 ));
    CascadeMux I__5152 (
            .O(N__29936),
            .I(N__29932));
    InMux I__5151 (
            .O(N__29935),
            .I(N__29928));
    InMux I__5150 (
            .O(N__29932),
            .I(N__29925));
    InMux I__5149 (
            .O(N__29931),
            .I(N__29922));
    LocalMux I__5148 (
            .O(N__29928),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    LocalMux I__5147 (
            .O(N__29925),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    LocalMux I__5146 (
            .O(N__29922),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    CascadeMux I__5145 (
            .O(N__29915),
            .I(N__29911));
    InMux I__5144 (
            .O(N__29914),
            .I(N__29905));
    InMux I__5143 (
            .O(N__29911),
            .I(N__29902));
    InMux I__5142 (
            .O(N__29910),
            .I(N__29899));
    InMux I__5141 (
            .O(N__29909),
            .I(N__29896));
    InMux I__5140 (
            .O(N__29908),
            .I(N__29893));
    LocalMux I__5139 (
            .O(N__29905),
            .I(N__29890));
    LocalMux I__5138 (
            .O(N__29902),
            .I(N__29885));
    LocalMux I__5137 (
            .O(N__29899),
            .I(N__29885));
    LocalMux I__5136 (
            .O(N__29896),
            .I(N__29880));
    LocalMux I__5135 (
            .O(N__29893),
            .I(N__29880));
    Span4Mux_v I__5134 (
            .O(N__29890),
            .I(N__29875));
    Span4Mux_v I__5133 (
            .O(N__29885),
            .I(N__29875));
    Span4Mux_v I__5132 (
            .O(N__29880),
            .I(N__29872));
    Odrv4 I__5131 (
            .O(N__29875),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__5130 (
            .O(N__29872),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__5129 (
            .O(N__29867),
            .I(N__29864));
    InMux I__5128 (
            .O(N__29864),
            .I(N__29861));
    LocalMux I__5127 (
            .O(N__29861),
            .I(N__29858));
    Span4Mux_h I__5126 (
            .O(N__29858),
            .I(N__29855));
    Odrv4 I__5125 (
            .O(N__29855),
            .I(\current_shift_inst.PI_CTRL.integrator_i_13 ));
    InMux I__5124 (
            .O(N__29852),
            .I(N__29849));
    LocalMux I__5123 (
            .O(N__29849),
            .I(N__29846));
    Span4Mux_h I__5122 (
            .O(N__29846),
            .I(N__29843));
    Odrv4 I__5121 (
            .O(N__29843),
            .I(\current_shift_inst.PI_CTRL.integrator_i_23 ));
    CascadeMux I__5120 (
            .O(N__29840),
            .I(N__29836));
    InMux I__5119 (
            .O(N__29839),
            .I(N__29831));
    InMux I__5118 (
            .O(N__29836),
            .I(N__29828));
    CascadeMux I__5117 (
            .O(N__29835),
            .I(N__29825));
    CascadeMux I__5116 (
            .O(N__29834),
            .I(N__29821));
    LocalMux I__5115 (
            .O(N__29831),
            .I(N__29818));
    LocalMux I__5114 (
            .O(N__29828),
            .I(N__29815));
    InMux I__5113 (
            .O(N__29825),
            .I(N__29812));
    InMux I__5112 (
            .O(N__29824),
            .I(N__29809));
    InMux I__5111 (
            .O(N__29821),
            .I(N__29806));
    Span4Mux_v I__5110 (
            .O(N__29818),
            .I(N__29801));
    Span4Mux_v I__5109 (
            .O(N__29815),
            .I(N__29801));
    LocalMux I__5108 (
            .O(N__29812),
            .I(N__29798));
    LocalMux I__5107 (
            .O(N__29809),
            .I(N__29795));
    LocalMux I__5106 (
            .O(N__29806),
            .I(N__29792));
    Span4Mux_h I__5105 (
            .O(N__29801),
            .I(N__29789));
    Span4Mux_h I__5104 (
            .O(N__29798),
            .I(N__29784));
    Span4Mux_h I__5103 (
            .O(N__29795),
            .I(N__29784));
    Odrv12 I__5102 (
            .O(N__29792),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__5101 (
            .O(N__29789),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__5100 (
            .O(N__29784),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__5099 (
            .O(N__29777),
            .I(N__29774));
    LocalMux I__5098 (
            .O(N__29774),
            .I(N__29771));
    Odrv12 I__5097 (
            .O(N__29771),
            .I(\current_shift_inst.PI_CTRL.integrator_i_16 ));
    InMux I__5096 (
            .O(N__29768),
            .I(N__29763));
    InMux I__5095 (
            .O(N__29767),
            .I(N__29760));
    InMux I__5094 (
            .O(N__29766),
            .I(N__29757));
    LocalMux I__5093 (
            .O(N__29763),
            .I(N__29752));
    LocalMux I__5092 (
            .O(N__29760),
            .I(N__29749));
    LocalMux I__5091 (
            .O(N__29757),
            .I(N__29746));
    InMux I__5090 (
            .O(N__29756),
            .I(N__29743));
    InMux I__5089 (
            .O(N__29755),
            .I(N__29740));
    Span4Mux_v I__5088 (
            .O(N__29752),
            .I(N__29737));
    Span4Mux_h I__5087 (
            .O(N__29749),
            .I(N__29734));
    Span4Mux_v I__5086 (
            .O(N__29746),
            .I(N__29729));
    LocalMux I__5085 (
            .O(N__29743),
            .I(N__29729));
    LocalMux I__5084 (
            .O(N__29740),
            .I(N__29726));
    Odrv4 I__5083 (
            .O(N__29737),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__5082 (
            .O(N__29734),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__5081 (
            .O(N__29729),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv12 I__5080 (
            .O(N__29726),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__5079 (
            .O(N__29717),
            .I(N__29714));
    LocalMux I__5078 (
            .O(N__29714),
            .I(N__29711));
    Odrv4 I__5077 (
            .O(N__29711),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ));
    CascadeMux I__5076 (
            .O(N__29708),
            .I(N__29705));
    InMux I__5075 (
            .O(N__29705),
            .I(N__29702));
    LocalMux I__5074 (
            .O(N__29702),
            .I(N__29699));
    Odrv12 I__5073 (
            .O(N__29699),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0 ));
    InMux I__5072 (
            .O(N__29696),
            .I(N__29693));
    LocalMux I__5071 (
            .O(N__29693),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ));
    InMux I__5070 (
            .O(N__29690),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ));
    InMux I__5069 (
            .O(N__29687),
            .I(N__29684));
    LocalMux I__5068 (
            .O(N__29684),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ));
    InMux I__5067 (
            .O(N__29681),
            .I(bfn_10_17_0_));
    InMux I__5066 (
            .O(N__29678),
            .I(N__29675));
    LocalMux I__5065 (
            .O(N__29675),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ));
    InMux I__5064 (
            .O(N__29672),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ));
    InMux I__5063 (
            .O(N__29669),
            .I(N__29666));
    LocalMux I__5062 (
            .O(N__29666),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ));
    InMux I__5061 (
            .O(N__29663),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ));
    InMux I__5060 (
            .O(N__29660),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ));
    InMux I__5059 (
            .O(N__29657),
            .I(N__29654));
    LocalMux I__5058 (
            .O(N__29654),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ));
    InMux I__5057 (
            .O(N__29651),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ));
    InMux I__5056 (
            .O(N__29648),
            .I(N__29645));
    LocalMux I__5055 (
            .O(N__29645),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ));
    InMux I__5054 (
            .O(N__29642),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ));
    InMux I__5053 (
            .O(N__29639),
            .I(N__29636));
    LocalMux I__5052 (
            .O(N__29636),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ));
    InMux I__5051 (
            .O(N__29633),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ));
    InMux I__5050 (
            .O(N__29630),
            .I(N__29627));
    LocalMux I__5049 (
            .O(N__29627),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ));
    InMux I__5048 (
            .O(N__29624),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ));
    InMux I__5047 (
            .O(N__29621),
            .I(N__29618));
    LocalMux I__5046 (
            .O(N__29618),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ));
    InMux I__5045 (
            .O(N__29615),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ));
    InMux I__5044 (
            .O(N__29612),
            .I(N__29609));
    LocalMux I__5043 (
            .O(N__29609),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ));
    InMux I__5042 (
            .O(N__29606),
            .I(bfn_10_16_0_));
    InMux I__5041 (
            .O(N__29603),
            .I(N__29600));
    LocalMux I__5040 (
            .O(N__29600),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ));
    InMux I__5039 (
            .O(N__29597),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ));
    InMux I__5038 (
            .O(N__29594),
            .I(N__29591));
    LocalMux I__5037 (
            .O(N__29591),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ));
    InMux I__5036 (
            .O(N__29588),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ));
    InMux I__5035 (
            .O(N__29585),
            .I(N__29582));
    LocalMux I__5034 (
            .O(N__29582),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ));
    InMux I__5033 (
            .O(N__29579),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ));
    CascadeMux I__5032 (
            .O(N__29576),
            .I(N__29573));
    InMux I__5031 (
            .O(N__29573),
            .I(N__29570));
    LocalMux I__5030 (
            .O(N__29570),
            .I(N__29567));
    Odrv4 I__5029 (
            .O(N__29567),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ));
    InMux I__5028 (
            .O(N__29564),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ));
    InMux I__5027 (
            .O(N__29561),
            .I(N__29558));
    LocalMux I__5026 (
            .O(N__29558),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ));
    InMux I__5025 (
            .O(N__29555),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ));
    InMux I__5024 (
            .O(N__29552),
            .I(N__29549));
    LocalMux I__5023 (
            .O(N__29549),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ));
    InMux I__5022 (
            .O(N__29546),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ));
    InMux I__5021 (
            .O(N__29543),
            .I(N__29540));
    LocalMux I__5020 (
            .O(N__29540),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_6 ));
    InMux I__5019 (
            .O(N__29537),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ));
    InMux I__5018 (
            .O(N__29534),
            .I(N__29531));
    LocalMux I__5017 (
            .O(N__29531),
            .I(N__29528));
    Odrv4 I__5016 (
            .O(N__29528),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_7 ));
    InMux I__5015 (
            .O(N__29525),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ));
    CascadeMux I__5014 (
            .O(N__29522),
            .I(N__29519));
    InMux I__5013 (
            .O(N__29519),
            .I(N__29516));
    LocalMux I__5012 (
            .O(N__29516),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_8 ));
    InMux I__5011 (
            .O(N__29513),
            .I(bfn_10_15_0_));
    InMux I__5010 (
            .O(N__29510),
            .I(N__29507));
    LocalMux I__5009 (
            .O(N__29507),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_9 ));
    InMux I__5008 (
            .O(N__29504),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ));
    InMux I__5007 (
            .O(N__29501),
            .I(N__29498));
    LocalMux I__5006 (
            .O(N__29498),
            .I(N__29495));
    Span4Mux_v I__5005 (
            .O(N__29495),
            .I(N__29492));
    Odrv4 I__5004 (
            .O(N__29492),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_10 ));
    InMux I__5003 (
            .O(N__29489),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ));
    InMux I__5002 (
            .O(N__29486),
            .I(N__29483));
    LocalMux I__5001 (
            .O(N__29483),
            .I(N__29480));
    Span4Mux_h I__5000 (
            .O(N__29480),
            .I(N__29477));
    Odrv4 I__4999 (
            .O(N__29477),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_11 ));
    InMux I__4998 (
            .O(N__29474),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ));
    InMux I__4997 (
            .O(N__29471),
            .I(N__29468));
    LocalMux I__4996 (
            .O(N__29468),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    InMux I__4995 (
            .O(N__29465),
            .I(N__29462));
    LocalMux I__4994 (
            .O(N__29462),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_12 ));
    InMux I__4993 (
            .O(N__29459),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ));
    InMux I__4992 (
            .O(N__29456),
            .I(N__29453));
    LocalMux I__4991 (
            .O(N__29453),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_13 ));
    InMux I__4990 (
            .O(N__29450),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ));
    InMux I__4989 (
            .O(N__29447),
            .I(N__29440));
    InMux I__4988 (
            .O(N__29446),
            .I(N__29440));
    InMux I__4987 (
            .O(N__29445),
            .I(N__29437));
    LocalMux I__4986 (
            .O(N__29440),
            .I(N__29434));
    LocalMux I__4985 (
            .O(N__29437),
            .I(N__29428));
    Span4Mux_h I__4984 (
            .O(N__29434),
            .I(N__29428));
    InMux I__4983 (
            .O(N__29433),
            .I(N__29425));
    Odrv4 I__4982 (
            .O(N__29428),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    LocalMux I__4981 (
            .O(N__29425),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__4980 (
            .O(N__29420),
            .I(N__29417));
    LocalMux I__4979 (
            .O(N__29417),
            .I(N__29413));
    InMux I__4978 (
            .O(N__29416),
            .I(N__29410));
    Odrv4 I__4977 (
            .O(N__29413),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    LocalMux I__4976 (
            .O(N__29410),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    InMux I__4975 (
            .O(N__29405),
            .I(N__29401));
    InMux I__4974 (
            .O(N__29404),
            .I(N__29398));
    LocalMux I__4973 (
            .O(N__29401),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    LocalMux I__4972 (
            .O(N__29398),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    InMux I__4971 (
            .O(N__29393),
            .I(N__29389));
    InMux I__4970 (
            .O(N__29392),
            .I(N__29386));
    LocalMux I__4969 (
            .O(N__29389),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    LocalMux I__4968 (
            .O(N__29386),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    InMux I__4967 (
            .O(N__29381),
            .I(N__29378));
    LocalMux I__4966 (
            .O(N__29378),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ));
    InMux I__4965 (
            .O(N__29375),
            .I(N__29372));
    LocalMux I__4964 (
            .O(N__29372),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ));
    InMux I__4963 (
            .O(N__29369),
            .I(N__29366));
    LocalMux I__4962 (
            .O(N__29366),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ));
    InMux I__4961 (
            .O(N__29363),
            .I(N__29360));
    LocalMux I__4960 (
            .O(N__29360),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ));
    InMux I__4959 (
            .O(N__29357),
            .I(N__29354));
    LocalMux I__4958 (
            .O(N__29354),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ));
    InMux I__4957 (
            .O(N__29351),
            .I(N__29348));
    LocalMux I__4956 (
            .O(N__29348),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_4 ));
    InMux I__4955 (
            .O(N__29345),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ));
    CascadeMux I__4954 (
            .O(N__29342),
            .I(N__29339));
    InMux I__4953 (
            .O(N__29339),
            .I(N__29336));
    LocalMux I__4952 (
            .O(N__29336),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_5 ));
    InMux I__4951 (
            .O(N__29333),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ));
    InMux I__4950 (
            .O(N__29330),
            .I(N__29327));
    LocalMux I__4949 (
            .O(N__29327),
            .I(N__29322));
    InMux I__4948 (
            .O(N__29326),
            .I(N__29319));
    InMux I__4947 (
            .O(N__29325),
            .I(N__29316));
    Span12Mux_h I__4946 (
            .O(N__29322),
            .I(N__29313));
    LocalMux I__4945 (
            .O(N__29319),
            .I(N__29310));
    LocalMux I__4944 (
            .O(N__29316),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv12 I__4943 (
            .O(N__29313),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv4 I__4942 (
            .O(N__29310),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__4941 (
            .O(N__29303),
            .I(N__29300));
    LocalMux I__4940 (
            .O(N__29300),
            .I(N__29297));
    Span4Mux_h I__4939 (
            .O(N__29297),
            .I(N__29293));
    InMux I__4938 (
            .O(N__29296),
            .I(N__29290));
    Span4Mux_v I__4937 (
            .O(N__29293),
            .I(N__29285));
    LocalMux I__4936 (
            .O(N__29290),
            .I(N__29282));
    InMux I__4935 (
            .O(N__29289),
            .I(N__29277));
    InMux I__4934 (
            .O(N__29288),
            .I(N__29277));
    Odrv4 I__4933 (
            .O(N__29285),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    Odrv4 I__4932 (
            .O(N__29282),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__4931 (
            .O(N__29277),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__4930 (
            .O(N__29270),
            .I(N__29267));
    LocalMux I__4929 (
            .O(N__29267),
            .I(N__29262));
    InMux I__4928 (
            .O(N__29266),
            .I(N__29259));
    InMux I__4927 (
            .O(N__29265),
            .I(N__29256));
    Span12Mux_v I__4926 (
            .O(N__29262),
            .I(N__29253));
    LocalMux I__4925 (
            .O(N__29259),
            .I(N__29250));
    LocalMux I__4924 (
            .O(N__29256),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    Odrv12 I__4923 (
            .O(N__29253),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    Odrv4 I__4922 (
            .O(N__29250),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__4921 (
            .O(N__29243),
            .I(N__29240));
    LocalMux I__4920 (
            .O(N__29240),
            .I(N__29237));
    Span4Mux_v I__4919 (
            .O(N__29237),
            .I(N__29231));
    InMux I__4918 (
            .O(N__29236),
            .I(N__29228));
    InMux I__4917 (
            .O(N__29235),
            .I(N__29223));
    InMux I__4916 (
            .O(N__29234),
            .I(N__29223));
    Odrv4 I__4915 (
            .O(N__29231),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__4914 (
            .O(N__29228),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__4913 (
            .O(N__29223),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__4912 (
            .O(N__29216),
            .I(N__29213));
    LocalMux I__4911 (
            .O(N__29213),
            .I(N__29210));
    Span4Mux_h I__4910 (
            .O(N__29210),
            .I(N__29206));
    InMux I__4909 (
            .O(N__29209),
            .I(N__29202));
    Span4Mux_v I__4908 (
            .O(N__29206),
            .I(N__29199));
    InMux I__4907 (
            .O(N__29205),
            .I(N__29196));
    LocalMux I__4906 (
            .O(N__29202),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    Odrv4 I__4905 (
            .O(N__29199),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    LocalMux I__4904 (
            .O(N__29196),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    InMux I__4903 (
            .O(N__29189),
            .I(N__29185));
    InMux I__4902 (
            .O(N__29188),
            .I(N__29181));
    LocalMux I__4901 (
            .O(N__29185),
            .I(N__29178));
    CascadeMux I__4900 (
            .O(N__29184),
            .I(N__29174));
    LocalMux I__4899 (
            .O(N__29181),
            .I(N__29171));
    Span4Mux_v I__4898 (
            .O(N__29178),
            .I(N__29168));
    InMux I__4897 (
            .O(N__29177),
            .I(N__29163));
    InMux I__4896 (
            .O(N__29174),
            .I(N__29163));
    Odrv4 I__4895 (
            .O(N__29171),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv4 I__4894 (
            .O(N__29168),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__4893 (
            .O(N__29163),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__4892 (
            .O(N__29156),
            .I(N__29153));
    LocalMux I__4891 (
            .O(N__29153),
            .I(N__29149));
    InMux I__4890 (
            .O(N__29152),
            .I(N__29146));
    Odrv4 I__4889 (
            .O(N__29149),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    LocalMux I__4888 (
            .O(N__29146),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    InMux I__4887 (
            .O(N__29141),
            .I(N__29136));
    InMux I__4886 (
            .O(N__29140),
            .I(N__29131));
    InMux I__4885 (
            .O(N__29139),
            .I(N__29131));
    LocalMux I__4884 (
            .O(N__29136),
            .I(N__29128));
    LocalMux I__4883 (
            .O(N__29131),
            .I(N__29125));
    Span4Mux_h I__4882 (
            .O(N__29128),
            .I(N__29121));
    Span4Mux_v I__4881 (
            .O(N__29125),
            .I(N__29118));
    InMux I__4880 (
            .O(N__29124),
            .I(N__29115));
    Odrv4 I__4879 (
            .O(N__29121),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__4878 (
            .O(N__29118),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__4877 (
            .O(N__29115),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    CascadeMux I__4876 (
            .O(N__29108),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_));
    CascadeMux I__4875 (
            .O(N__29105),
            .I(N__29102));
    InMux I__4874 (
            .O(N__29102),
            .I(N__29096));
    InMux I__4873 (
            .O(N__29101),
            .I(N__29096));
    LocalMux I__4872 (
            .O(N__29096),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ));
    InMux I__4871 (
            .O(N__29093),
            .I(N__29090));
    LocalMux I__4870 (
            .O(N__29090),
            .I(N__29087));
    Span4Mux_h I__4869 (
            .O(N__29087),
            .I(N__29083));
    InMux I__4868 (
            .O(N__29086),
            .I(N__29080));
    Odrv4 I__4867 (
            .O(N__29083),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    LocalMux I__4866 (
            .O(N__29080),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__4865 (
            .O(N__29075),
            .I(N__29068));
    InMux I__4864 (
            .O(N__29074),
            .I(N__29068));
    InMux I__4863 (
            .O(N__29073),
            .I(N__29064));
    LocalMux I__4862 (
            .O(N__29068),
            .I(N__29061));
    InMux I__4861 (
            .O(N__29067),
            .I(N__29058));
    LocalMux I__4860 (
            .O(N__29064),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv4 I__4859 (
            .O(N__29061),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__4858 (
            .O(N__29058),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    CascadeMux I__4857 (
            .O(N__29051),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24_cascade_));
    CascadeMux I__4856 (
            .O(N__29048),
            .I(N__29045));
    InMux I__4855 (
            .O(N__29045),
            .I(N__29041));
    InMux I__4854 (
            .O(N__29044),
            .I(N__29038));
    LocalMux I__4853 (
            .O(N__29041),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    LocalMux I__4852 (
            .O(N__29038),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    InMux I__4851 (
            .O(N__29033),
            .I(N__29030));
    LocalMux I__4850 (
            .O(N__29030),
            .I(N__29027));
    Span4Mux_v I__4849 (
            .O(N__29027),
            .I(N__29023));
    InMux I__4848 (
            .O(N__29026),
            .I(N__29020));
    Odrv4 I__4847 (
            .O(N__29023),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    LocalMux I__4846 (
            .O(N__29020),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    CascadeMux I__4845 (
            .O(N__29015),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_));
    InMux I__4844 (
            .O(N__29012),
            .I(N__29009));
    LocalMux I__4843 (
            .O(N__29009),
            .I(N__29006));
    Span4Mux_h I__4842 (
            .O(N__29006),
            .I(N__29000));
    InMux I__4841 (
            .O(N__29005),
            .I(N__28995));
    InMux I__4840 (
            .O(N__29004),
            .I(N__28995));
    InMux I__4839 (
            .O(N__29003),
            .I(N__28992));
    Odrv4 I__4838 (
            .O(N__29000),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    LocalMux I__4837 (
            .O(N__28995),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    LocalMux I__4836 (
            .O(N__28992),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    CascadeMux I__4835 (
            .O(N__28985),
            .I(N__28982));
    InMux I__4834 (
            .O(N__28982),
            .I(N__28976));
    InMux I__4833 (
            .O(N__28981),
            .I(N__28976));
    LocalMux I__4832 (
            .O(N__28976),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__4831 (
            .O(N__28973),
            .I(N__28970));
    LocalMux I__4830 (
            .O(N__28970),
            .I(N__28967));
    Span4Mux_h I__4829 (
            .O(N__28967),
            .I(N__28963));
    InMux I__4828 (
            .O(N__28966),
            .I(N__28960));
    Odrv4 I__4827 (
            .O(N__28963),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    LocalMux I__4826 (
            .O(N__28960),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    CascadeMux I__4825 (
            .O(N__28955),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_));
    InMux I__4824 (
            .O(N__28952),
            .I(N__28949));
    LocalMux I__4823 (
            .O(N__28949),
            .I(N__28944));
    InMux I__4822 (
            .O(N__28948),
            .I(N__28939));
    InMux I__4821 (
            .O(N__28947),
            .I(N__28939));
    Span4Mux_h I__4820 (
            .O(N__28944),
            .I(N__28933));
    LocalMux I__4819 (
            .O(N__28939),
            .I(N__28933));
    InMux I__4818 (
            .O(N__28938),
            .I(N__28930));
    Odrv4 I__4817 (
            .O(N__28933),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__4816 (
            .O(N__28930),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__4815 (
            .O(N__28925),
            .I(N__28919));
    InMux I__4814 (
            .O(N__28924),
            .I(N__28919));
    LocalMux I__4813 (
            .O(N__28919),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__4812 (
            .O(N__28916),
            .I(N__28913));
    LocalMux I__4811 (
            .O(N__28913),
            .I(N__28910));
    Span4Mux_h I__4810 (
            .O(N__28910),
            .I(N__28906));
    InMux I__4809 (
            .O(N__28909),
            .I(N__28903));
    Odrv4 I__4808 (
            .O(N__28906),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    LocalMux I__4807 (
            .O(N__28903),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    CascadeMux I__4806 (
            .O(N__28898),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_));
    InMux I__4805 (
            .O(N__28895),
            .I(N__28890));
    InMux I__4804 (
            .O(N__28894),
            .I(N__28885));
    InMux I__4803 (
            .O(N__28893),
            .I(N__28885));
    LocalMux I__4802 (
            .O(N__28890),
            .I(N__28881));
    LocalMux I__4801 (
            .O(N__28885),
            .I(N__28878));
    InMux I__4800 (
            .O(N__28884),
            .I(N__28875));
    Odrv4 I__4799 (
            .O(N__28881),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv4 I__4798 (
            .O(N__28878),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__4797 (
            .O(N__28875),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__4796 (
            .O(N__28868),
            .I(N__28862));
    InMux I__4795 (
            .O(N__28867),
            .I(N__28862));
    LocalMux I__4794 (
            .O(N__28862),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    InMux I__4793 (
            .O(N__28859),
            .I(N__28856));
    LocalMux I__4792 (
            .O(N__28856),
            .I(N__28853));
    Span4Mux_v I__4791 (
            .O(N__28853),
            .I(N__28848));
    InMux I__4790 (
            .O(N__28852),
            .I(N__28845));
    InMux I__4789 (
            .O(N__28851),
            .I(N__28842));
    Span4Mux_v I__4788 (
            .O(N__28848),
            .I(N__28839));
    LocalMux I__4787 (
            .O(N__28845),
            .I(N__28836));
    LocalMux I__4786 (
            .O(N__28842),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__4785 (
            .O(N__28839),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__4784 (
            .O(N__28836),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__4783 (
            .O(N__28829),
            .I(N__28826));
    LocalMux I__4782 (
            .O(N__28826),
            .I(N__28823));
    Span4Mux_h I__4781 (
            .O(N__28823),
            .I(N__28819));
    InMux I__4780 (
            .O(N__28822),
            .I(N__28816));
    Span4Mux_v I__4779 (
            .O(N__28819),
            .I(N__28811));
    LocalMux I__4778 (
            .O(N__28816),
            .I(N__28808));
    InMux I__4777 (
            .O(N__28815),
            .I(N__28803));
    InMux I__4776 (
            .O(N__28814),
            .I(N__28803));
    Odrv4 I__4775 (
            .O(N__28811),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    Odrv4 I__4774 (
            .O(N__28808),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__4773 (
            .O(N__28803),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    CascadeMux I__4772 (
            .O(N__28796),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_));
    InMux I__4771 (
            .O(N__28793),
            .I(N__28787));
    InMux I__4770 (
            .O(N__28792),
            .I(N__28784));
    InMux I__4769 (
            .O(N__28791),
            .I(N__28779));
    InMux I__4768 (
            .O(N__28790),
            .I(N__28779));
    LocalMux I__4767 (
            .O(N__28787),
            .I(N__28776));
    LocalMux I__4766 (
            .O(N__28784),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    LocalMux I__4765 (
            .O(N__28779),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__4764 (
            .O(N__28776),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__4763 (
            .O(N__28769),
            .I(N__28765));
    CascadeMux I__4762 (
            .O(N__28768),
            .I(N__28762));
    LocalMux I__4761 (
            .O(N__28765),
            .I(N__28759));
    InMux I__4760 (
            .O(N__28762),
            .I(N__28756));
    Odrv4 I__4759 (
            .O(N__28759),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    LocalMux I__4758 (
            .O(N__28756),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    CascadeMux I__4757 (
            .O(N__28751),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31_cascade_));
    InMux I__4756 (
            .O(N__28748),
            .I(N__28745));
    LocalMux I__4755 (
            .O(N__28745),
            .I(N__28739));
    InMux I__4754 (
            .O(N__28744),
            .I(N__28736));
    InMux I__4753 (
            .O(N__28743),
            .I(N__28731));
    InMux I__4752 (
            .O(N__28742),
            .I(N__28731));
    Span4Mux_h I__4751 (
            .O(N__28739),
            .I(N__28728));
    LocalMux I__4750 (
            .O(N__28736),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    LocalMux I__4749 (
            .O(N__28731),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__4748 (
            .O(N__28728),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    CascadeMux I__4747 (
            .O(N__28721),
            .I(N__28716));
    CascadeMux I__4746 (
            .O(N__28720),
            .I(N__28713));
    InMux I__4745 (
            .O(N__28719),
            .I(N__28706));
    InMux I__4744 (
            .O(N__28716),
            .I(N__28706));
    InMux I__4743 (
            .O(N__28713),
            .I(N__28706));
    LocalMux I__4742 (
            .O(N__28706),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    InMux I__4741 (
            .O(N__28703),
            .I(N__28694));
    InMux I__4740 (
            .O(N__28702),
            .I(N__28694));
    InMux I__4739 (
            .O(N__28701),
            .I(N__28694));
    LocalMux I__4738 (
            .O(N__28694),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    InMux I__4737 (
            .O(N__28691),
            .I(N__28688));
    LocalMux I__4736 (
            .O(N__28688),
            .I(N__28684));
    InMux I__4735 (
            .O(N__28687),
            .I(N__28681));
    Odrv4 I__4734 (
            .O(N__28684),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    LocalMux I__4733 (
            .O(N__28681),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    InMux I__4732 (
            .O(N__28676),
            .I(N__28670));
    InMux I__4731 (
            .O(N__28675),
            .I(N__28665));
    InMux I__4730 (
            .O(N__28674),
            .I(N__28665));
    InMux I__4729 (
            .O(N__28673),
            .I(N__28662));
    LocalMux I__4728 (
            .O(N__28670),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__4727 (
            .O(N__28665),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__4726 (
            .O(N__28662),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__4725 (
            .O(N__28655),
            .I(N__28651));
    InMux I__4724 (
            .O(N__28654),
            .I(N__28646));
    LocalMux I__4723 (
            .O(N__28651),
            .I(N__28643));
    InMux I__4722 (
            .O(N__28650),
            .I(N__28638));
    InMux I__4721 (
            .O(N__28649),
            .I(N__28638));
    LocalMux I__4720 (
            .O(N__28646),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    Odrv4 I__4719 (
            .O(N__28643),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    LocalMux I__4718 (
            .O(N__28638),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__4717 (
            .O(N__28631),
            .I(N__28626));
    InMux I__4716 (
            .O(N__28630),
            .I(N__28623));
    InMux I__4715 (
            .O(N__28629),
            .I(N__28620));
    LocalMux I__4714 (
            .O(N__28626),
            .I(N__28617));
    LocalMux I__4713 (
            .O(N__28623),
            .I(N__28614));
    LocalMux I__4712 (
            .O(N__28620),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv4 I__4711 (
            .O(N__28617),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv12 I__4710 (
            .O(N__28614),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    InMux I__4709 (
            .O(N__28607),
            .I(N__28599));
    InMux I__4708 (
            .O(N__28606),
            .I(N__28599));
    CascadeMux I__4707 (
            .O(N__28605),
            .I(N__28596));
    InMux I__4706 (
            .O(N__28604),
            .I(N__28593));
    LocalMux I__4705 (
            .O(N__28599),
            .I(N__28590));
    InMux I__4704 (
            .O(N__28596),
            .I(N__28587));
    LocalMux I__4703 (
            .O(N__28593),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__4702 (
            .O(N__28590),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    LocalMux I__4701 (
            .O(N__28587),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__4700 (
            .O(N__28580),
            .I(N__28577));
    LocalMux I__4699 (
            .O(N__28577),
            .I(N__28574));
    Span4Mux_v I__4698 (
            .O(N__28574),
            .I(N__28570));
    InMux I__4697 (
            .O(N__28573),
            .I(N__28567));
    Odrv4 I__4696 (
            .O(N__28570),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__4695 (
            .O(N__28567),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    InMux I__4694 (
            .O(N__28562),
            .I(N__28559));
    LocalMux I__4693 (
            .O(N__28559),
            .I(N__28554));
    InMux I__4692 (
            .O(N__28558),
            .I(N__28551));
    CascadeMux I__4691 (
            .O(N__28557),
            .I(N__28548));
    Span4Mux_v I__4690 (
            .O(N__28554),
            .I(N__28542));
    LocalMux I__4689 (
            .O(N__28551),
            .I(N__28542));
    InMux I__4688 (
            .O(N__28548),
            .I(N__28539));
    InMux I__4687 (
            .O(N__28547),
            .I(N__28536));
    Span4Mux_h I__4686 (
            .O(N__28542),
            .I(N__28533));
    LocalMux I__4685 (
            .O(N__28539),
            .I(N__28530));
    LocalMux I__4684 (
            .O(N__28536),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__4683 (
            .O(N__28533),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__4682 (
            .O(N__28530),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    CascadeMux I__4681 (
            .O(N__28523),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_ ));
    InMux I__4680 (
            .O(N__28520),
            .I(N__28517));
    LocalMux I__4679 (
            .O(N__28517),
            .I(N__28514));
    Odrv4 I__4678 (
            .O(N__28514),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    InMux I__4677 (
            .O(N__28511),
            .I(N__28508));
    LocalMux I__4676 (
            .O(N__28508),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    InMux I__4675 (
            .O(N__28505),
            .I(N__28502));
    LocalMux I__4674 (
            .O(N__28502),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    InMux I__4673 (
            .O(N__28499),
            .I(N__28496));
    LocalMux I__4672 (
            .O(N__28496),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ));
    InMux I__4671 (
            .O(N__28493),
            .I(N__28490));
    LocalMux I__4670 (
            .O(N__28490),
            .I(N__28486));
    InMux I__4669 (
            .O(N__28489),
            .I(N__28483));
    Odrv4 I__4668 (
            .O(N__28486),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    LocalMux I__4667 (
            .O(N__28483),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    CascadeMux I__4666 (
            .O(N__28478),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ));
    InMux I__4665 (
            .O(N__28475),
            .I(N__28472));
    LocalMux I__4664 (
            .O(N__28472),
            .I(N__28469));
    Odrv12 I__4663 (
            .O(N__28469),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ));
    CascadeMux I__4662 (
            .O(N__28466),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ));
    InMux I__4661 (
            .O(N__28463),
            .I(N__28459));
    InMux I__4660 (
            .O(N__28462),
            .I(N__28456));
    LocalMux I__4659 (
            .O(N__28459),
            .I(N__28451));
    LocalMux I__4658 (
            .O(N__28456),
            .I(N__28448));
    InMux I__4657 (
            .O(N__28455),
            .I(N__28443));
    InMux I__4656 (
            .O(N__28454),
            .I(N__28443));
    Odrv4 I__4655 (
            .O(N__28451),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__4654 (
            .O(N__28448),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    LocalMux I__4653 (
            .O(N__28443),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    CascadeMux I__4652 (
            .O(N__28436),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__4651 (
            .O(N__28433),
            .I(N__28430));
    LocalMux I__4650 (
            .O(N__28430),
            .I(N__28426));
    InMux I__4649 (
            .O(N__28429),
            .I(N__28423));
    Span4Mux_v I__4648 (
            .O(N__28426),
            .I(N__28417));
    LocalMux I__4647 (
            .O(N__28423),
            .I(N__28417));
    InMux I__4646 (
            .O(N__28422),
            .I(N__28414));
    Span4Mux_h I__4645 (
            .O(N__28417),
            .I(N__28411));
    LocalMux I__4644 (
            .O(N__28414),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    Odrv4 I__4643 (
            .O(N__28411),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    InMux I__4642 (
            .O(N__28406),
            .I(N__28403));
    LocalMux I__4641 (
            .O(N__28403),
            .I(N__28400));
    Span4Mux_v I__4640 (
            .O(N__28400),
            .I(N__28396));
    InMux I__4639 (
            .O(N__28399),
            .I(N__28393));
    Odrv4 I__4638 (
            .O(N__28396),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__4637 (
            .O(N__28393),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    CascadeMux I__4636 (
            .O(N__28388),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_));
    InMux I__4635 (
            .O(N__28385),
            .I(N__28382));
    LocalMux I__4634 (
            .O(N__28382),
            .I(N__28376));
    InMux I__4633 (
            .O(N__28381),
            .I(N__28373));
    InMux I__4632 (
            .O(N__28380),
            .I(N__28368));
    InMux I__4631 (
            .O(N__28379),
            .I(N__28368));
    Odrv4 I__4630 (
            .O(N__28376),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__4629 (
            .O(N__28373),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__4628 (
            .O(N__28368),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__4627 (
            .O(N__28361),
            .I(N__28358));
    LocalMux I__4626 (
            .O(N__28358),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ));
    InMux I__4625 (
            .O(N__28355),
            .I(N__28352));
    LocalMux I__4624 (
            .O(N__28352),
            .I(N__28348));
    InMux I__4623 (
            .O(N__28351),
            .I(N__28345));
    Odrv4 I__4622 (
            .O(N__28348),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    LocalMux I__4621 (
            .O(N__28345),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    CascadeMux I__4620 (
            .O(N__28340),
            .I(elapsed_time_ns_1_RNILK91B_0_9_cascade_));
    InMux I__4619 (
            .O(N__28337),
            .I(N__28331));
    InMux I__4618 (
            .O(N__28336),
            .I(N__28324));
    InMux I__4617 (
            .O(N__28335),
            .I(N__28324));
    InMux I__4616 (
            .O(N__28334),
            .I(N__28324));
    LocalMux I__4615 (
            .O(N__28331),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    LocalMux I__4614 (
            .O(N__28324),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    CascadeMux I__4613 (
            .O(N__28319),
            .I(N__28316));
    InMux I__4612 (
            .O(N__28316),
            .I(N__28313));
    LocalMux I__4611 (
            .O(N__28313),
            .I(N__28310));
    Odrv4 I__4610 (
            .O(N__28310),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__4609 (
            .O(N__28307),
            .I(N__28304));
    LocalMux I__4608 (
            .O(N__28304),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__4607 (
            .O(N__28301),
            .I(N__28298));
    LocalMux I__4606 (
            .O(N__28298),
            .I(N__28294));
    CascadeMux I__4605 (
            .O(N__28297),
            .I(N__28289));
    Span4Mux_h I__4604 (
            .O(N__28294),
            .I(N__28286));
    InMux I__4603 (
            .O(N__28293),
            .I(N__28283));
    InMux I__4602 (
            .O(N__28292),
            .I(N__28280));
    InMux I__4601 (
            .O(N__28289),
            .I(N__28277));
    Span4Mux_v I__4600 (
            .O(N__28286),
            .I(N__28272));
    LocalMux I__4599 (
            .O(N__28283),
            .I(N__28272));
    LocalMux I__4598 (
            .O(N__28280),
            .I(N__28269));
    LocalMux I__4597 (
            .O(N__28277),
            .I(N__28264));
    Span4Mux_h I__4596 (
            .O(N__28272),
            .I(N__28264));
    Span4Mux_h I__4595 (
            .O(N__28269),
            .I(N__28261));
    Span4Mux_h I__4594 (
            .O(N__28264),
            .I(N__28258));
    Odrv4 I__4593 (
            .O(N__28261),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__4592 (
            .O(N__28258),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__4591 (
            .O(N__28253),
            .I(N__28250));
    InMux I__4590 (
            .O(N__28250),
            .I(N__28247));
    LocalMux I__4589 (
            .O(N__28247),
            .I(N__28244));
    Span4Mux_v I__4588 (
            .O(N__28244),
            .I(N__28241));
    Span4Mux_h I__4587 (
            .O(N__28241),
            .I(N__28238));
    Odrv4 I__4586 (
            .O(N__28238),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__4585 (
            .O(N__28235),
            .I(N__28230));
    InMux I__4584 (
            .O(N__28234),
            .I(N__28226));
    InMux I__4583 (
            .O(N__28233),
            .I(N__28223));
    InMux I__4582 (
            .O(N__28230),
            .I(N__28220));
    InMux I__4581 (
            .O(N__28229),
            .I(N__28217));
    LocalMux I__4580 (
            .O(N__28226),
            .I(N__28214));
    LocalMux I__4579 (
            .O(N__28223),
            .I(N__28209));
    LocalMux I__4578 (
            .O(N__28220),
            .I(N__28209));
    LocalMux I__4577 (
            .O(N__28217),
            .I(N__28206));
    Span4Mux_h I__4576 (
            .O(N__28214),
            .I(N__28200));
    Span4Mux_h I__4575 (
            .O(N__28209),
            .I(N__28200));
    Span4Mux_h I__4574 (
            .O(N__28206),
            .I(N__28197));
    InMux I__4573 (
            .O(N__28205),
            .I(N__28194));
    Odrv4 I__4572 (
            .O(N__28200),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__4571 (
            .O(N__28197),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__4570 (
            .O(N__28194),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__4569 (
            .O(N__28187),
            .I(N__28183));
    CascadeMux I__4568 (
            .O(N__28186),
            .I(N__28180));
    LocalMux I__4567 (
            .O(N__28183),
            .I(N__28176));
    InMux I__4566 (
            .O(N__28180),
            .I(N__28171));
    InMux I__4565 (
            .O(N__28179),
            .I(N__28171));
    Span4Mux_h I__4564 (
            .O(N__28176),
            .I(N__28166));
    LocalMux I__4563 (
            .O(N__28171),
            .I(N__28166));
    Span4Mux_v I__4562 (
            .O(N__28166),
            .I(N__28163));
    Span4Mux_v I__4561 (
            .O(N__28163),
            .I(N__28160));
    Span4Mux_v I__4560 (
            .O(N__28160),
            .I(N__28157));
    Odrv4 I__4559 (
            .O(N__28157),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__4558 (
            .O(N__28154),
            .I(N__28151));
    LocalMux I__4557 (
            .O(N__28151),
            .I(N__28147));
    InMux I__4556 (
            .O(N__28150),
            .I(N__28144));
    Span4Mux_h I__4555 (
            .O(N__28147),
            .I(N__28139));
    LocalMux I__4554 (
            .O(N__28144),
            .I(N__28139));
    Span4Mux_v I__4553 (
            .O(N__28139),
            .I(N__28136));
    Span4Mux_v I__4552 (
            .O(N__28136),
            .I(N__28131));
    InMux I__4551 (
            .O(N__28135),
            .I(N__28126));
    InMux I__4550 (
            .O(N__28134),
            .I(N__28126));
    Span4Mux_v I__4549 (
            .O(N__28131),
            .I(N__28123));
    LocalMux I__4548 (
            .O(N__28126),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__4547 (
            .O(N__28123),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__4546 (
            .O(N__28118),
            .I(N__28115));
    GlobalMux I__4545 (
            .O(N__28115),
            .I(N__28112));
    gio2CtrlBuf I__4544 (
            .O(N__28112),
            .I(delay_tr_input_c_g));
    IoInMux I__4543 (
            .O(N__28109),
            .I(N__28106));
    LocalMux I__4542 (
            .O(N__28106),
            .I(N__28103));
    Odrv12 I__4541 (
            .O(N__28103),
            .I(s3_phy_c));
    InMux I__4540 (
            .O(N__28100),
            .I(N__28097));
    LocalMux I__4539 (
            .O(N__28097),
            .I(N__28094));
    Glb2LocalMux I__4538 (
            .O(N__28094),
            .I(N__28091));
    GlobalMux I__4537 (
            .O(N__28091),
            .I(clk_12mhz));
    IoInMux I__4536 (
            .O(N__28088),
            .I(N__28085));
    LocalMux I__4535 (
            .O(N__28085),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__4534 (
            .O(N__28082),
            .I(N__28079));
    LocalMux I__4533 (
            .O(N__28079),
            .I(N__28076));
    Span4Mux_h I__4532 (
            .O(N__28076),
            .I(N__28073));
    Odrv4 I__4531 (
            .O(N__28073),
            .I(il_max_comp1_c));
    InMux I__4530 (
            .O(N__28070),
            .I(N__28067));
    LocalMux I__4529 (
            .O(N__28067),
            .I(\current_shift_inst.PI_CTRL.integrator_i_10 ));
    CascadeMux I__4528 (
            .O(N__28064),
            .I(N__28061));
    InMux I__4527 (
            .O(N__28061),
            .I(N__28057));
    CascadeMux I__4526 (
            .O(N__28060),
            .I(N__28054));
    LocalMux I__4525 (
            .O(N__28057),
            .I(N__28049));
    InMux I__4524 (
            .O(N__28054),
            .I(N__28044));
    InMux I__4523 (
            .O(N__28053),
            .I(N__28044));
    InMux I__4522 (
            .O(N__28052),
            .I(N__28040));
    Span4Mux_v I__4521 (
            .O(N__28049),
            .I(N__28035));
    LocalMux I__4520 (
            .O(N__28044),
            .I(N__28035));
    InMux I__4519 (
            .O(N__28043),
            .I(N__28032));
    LocalMux I__4518 (
            .O(N__28040),
            .I(N__28027));
    Span4Mux_h I__4517 (
            .O(N__28035),
            .I(N__28027));
    LocalMux I__4516 (
            .O(N__28032),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__4515 (
            .O(N__28027),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__4514 (
            .O(N__28022),
            .I(N__28019));
    InMux I__4513 (
            .O(N__28019),
            .I(N__28016));
    LocalMux I__4512 (
            .O(N__28016),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0 ));
    InMux I__4511 (
            .O(N__28013),
            .I(N__28008));
    InMux I__4510 (
            .O(N__28012),
            .I(N__28005));
    CascadeMux I__4509 (
            .O(N__28011),
            .I(N__28001));
    LocalMux I__4508 (
            .O(N__28008),
            .I(N__27998));
    LocalMux I__4507 (
            .O(N__28005),
            .I(N__27995));
    InMux I__4506 (
            .O(N__28004),
            .I(N__27991));
    InMux I__4505 (
            .O(N__28001),
            .I(N__27988));
    Span4Mux_v I__4504 (
            .O(N__27998),
            .I(N__27983));
    Span4Mux_v I__4503 (
            .O(N__27995),
            .I(N__27983));
    InMux I__4502 (
            .O(N__27994),
            .I(N__27980));
    LocalMux I__4501 (
            .O(N__27991),
            .I(N__27975));
    LocalMux I__4500 (
            .O(N__27988),
            .I(N__27975));
    Odrv4 I__4499 (
            .O(N__27983),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__4498 (
            .O(N__27980),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv12 I__4497 (
            .O(N__27975),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    CascadeMux I__4496 (
            .O(N__27968),
            .I(N__27965));
    InMux I__4495 (
            .O(N__27965),
            .I(N__27962));
    LocalMux I__4494 (
            .O(N__27962),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0 ));
    InMux I__4493 (
            .O(N__27959),
            .I(N__27956));
    LocalMux I__4492 (
            .O(N__27956),
            .I(N__27953));
    Odrv4 I__4491 (
            .O(N__27953),
            .I(\current_shift_inst.PI_CTRL.integrator_i_6 ));
    CascadeMux I__4490 (
            .O(N__27950),
            .I(N__27946));
    InMux I__4489 (
            .O(N__27949),
            .I(N__27943));
    InMux I__4488 (
            .O(N__27946),
            .I(N__27940));
    LocalMux I__4487 (
            .O(N__27943),
            .I(N__27935));
    LocalMux I__4486 (
            .O(N__27940),
            .I(N__27932));
    InMux I__4485 (
            .O(N__27939),
            .I(N__27926));
    InMux I__4484 (
            .O(N__27938),
            .I(N__27926));
    Span4Mux_h I__4483 (
            .O(N__27935),
            .I(N__27921));
    Span4Mux_h I__4482 (
            .O(N__27932),
            .I(N__27921));
    InMux I__4481 (
            .O(N__27931),
            .I(N__27918));
    LocalMux I__4480 (
            .O(N__27926),
            .I(N__27915));
    Odrv4 I__4479 (
            .O(N__27921),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__4478 (
            .O(N__27918),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__4477 (
            .O(N__27915),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    CascadeMux I__4476 (
            .O(N__27908),
            .I(N__27905));
    InMux I__4475 (
            .O(N__27905),
            .I(N__27902));
    LocalMux I__4474 (
            .O(N__27902),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0 ));
    CascadeMux I__4473 (
            .O(N__27899),
            .I(N__27896));
    InMux I__4472 (
            .O(N__27896),
            .I(N__27893));
    LocalMux I__4471 (
            .O(N__27893),
            .I(N__27890));
    Odrv4 I__4470 (
            .O(N__27890),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0 ));
    CascadeMux I__4469 (
            .O(N__27887),
            .I(N__27884));
    InMux I__4468 (
            .O(N__27884),
            .I(N__27881));
    LocalMux I__4467 (
            .O(N__27881),
            .I(N__27878));
    Odrv4 I__4466 (
            .O(N__27878),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10 ));
    InMux I__4465 (
            .O(N__27875),
            .I(N__27872));
    LocalMux I__4464 (
            .O(N__27872),
            .I(N__27869));
    Odrv4 I__4463 (
            .O(N__27869),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__4462 (
            .O(N__27866),
            .I(N__27863));
    InMux I__4461 (
            .O(N__27863),
            .I(N__27858));
    InMux I__4460 (
            .O(N__27862),
            .I(N__27855));
    InMux I__4459 (
            .O(N__27861),
            .I(N__27851));
    LocalMux I__4458 (
            .O(N__27858),
            .I(N__27846));
    LocalMux I__4457 (
            .O(N__27855),
            .I(N__27846));
    InMux I__4456 (
            .O(N__27854),
            .I(N__27843));
    LocalMux I__4455 (
            .O(N__27851),
            .I(N__27838));
    Span4Mux_h I__4454 (
            .O(N__27846),
            .I(N__27838));
    LocalMux I__4453 (
            .O(N__27843),
            .I(N__27832));
    Span4Mux_v I__4452 (
            .O(N__27838),
            .I(N__27832));
    InMux I__4451 (
            .O(N__27837),
            .I(N__27829));
    Odrv4 I__4450 (
            .O(N__27832),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__4449 (
            .O(N__27829),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__4448 (
            .O(N__27824),
            .I(N__27821));
    LocalMux I__4447 (
            .O(N__27821),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__4446 (
            .O(N__27818),
            .I(N__27814));
    CascadeMux I__4445 (
            .O(N__27817),
            .I(N__27810));
    LocalMux I__4444 (
            .O(N__27814),
            .I(N__27805));
    InMux I__4443 (
            .O(N__27813),
            .I(N__27802));
    InMux I__4442 (
            .O(N__27810),
            .I(N__27799));
    InMux I__4441 (
            .O(N__27809),
            .I(N__27796));
    InMux I__4440 (
            .O(N__27808),
            .I(N__27793));
    Span4Mux_v I__4439 (
            .O(N__27805),
            .I(N__27790));
    LocalMux I__4438 (
            .O(N__27802),
            .I(N__27783));
    LocalMux I__4437 (
            .O(N__27799),
            .I(N__27783));
    LocalMux I__4436 (
            .O(N__27796),
            .I(N__27783));
    LocalMux I__4435 (
            .O(N__27793),
            .I(N__27780));
    Span4Mux_v I__4434 (
            .O(N__27790),
            .I(N__27775));
    Span4Mux_v I__4433 (
            .O(N__27783),
            .I(N__27775));
    Span4Mux_h I__4432 (
            .O(N__27780),
            .I(N__27772));
    Odrv4 I__4431 (
            .O(N__27775),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__4430 (
            .O(N__27772),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__4429 (
            .O(N__27767),
            .I(N__27764));
    LocalMux I__4428 (
            .O(N__27764),
            .I(\current_shift_inst.PI_CTRL.integrator_i_14 ));
    CascadeMux I__4427 (
            .O(N__27761),
            .I(N__27758));
    InMux I__4426 (
            .O(N__27758),
            .I(N__27755));
    LocalMux I__4425 (
            .O(N__27755),
            .I(N__27752));
    Odrv4 I__4424 (
            .O(N__27752),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0 ));
    CascadeMux I__4423 (
            .O(N__27749),
            .I(N__27745));
    InMux I__4422 (
            .O(N__27748),
            .I(N__27740));
    InMux I__4421 (
            .O(N__27745),
            .I(N__27737));
    InMux I__4420 (
            .O(N__27744),
            .I(N__27734));
    InMux I__4419 (
            .O(N__27743),
            .I(N__27730));
    LocalMux I__4418 (
            .O(N__27740),
            .I(N__27727));
    LocalMux I__4417 (
            .O(N__27737),
            .I(N__27722));
    LocalMux I__4416 (
            .O(N__27734),
            .I(N__27722));
    InMux I__4415 (
            .O(N__27733),
            .I(N__27719));
    LocalMux I__4414 (
            .O(N__27730),
            .I(N__27716));
    Span12Mux_h I__4413 (
            .O(N__27727),
            .I(N__27709));
    Span12Mux_s7_h I__4412 (
            .O(N__27722),
            .I(N__27709));
    LocalMux I__4411 (
            .O(N__27719),
            .I(N__27709));
    Odrv12 I__4410 (
            .O(N__27716),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv12 I__4409 (
            .O(N__27709),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__4408 (
            .O(N__27704),
            .I(N__27701));
    InMux I__4407 (
            .O(N__27701),
            .I(N__27698));
    LocalMux I__4406 (
            .O(N__27698),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0 ));
    InMux I__4405 (
            .O(N__27695),
            .I(N__27689));
    InMux I__4404 (
            .O(N__27694),
            .I(N__27686));
    InMux I__4403 (
            .O(N__27693),
            .I(N__27680));
    InMux I__4402 (
            .O(N__27692),
            .I(N__27680));
    LocalMux I__4401 (
            .O(N__27689),
            .I(N__27677));
    LocalMux I__4400 (
            .O(N__27686),
            .I(N__27674));
    InMux I__4399 (
            .O(N__27685),
            .I(N__27671));
    LocalMux I__4398 (
            .O(N__27680),
            .I(N__27668));
    Span4Mux_h I__4397 (
            .O(N__27677),
            .I(N__27665));
    Span4Mux_h I__4396 (
            .O(N__27674),
            .I(N__27658));
    LocalMux I__4395 (
            .O(N__27671),
            .I(N__27658));
    Span4Mux_h I__4394 (
            .O(N__27668),
            .I(N__27658));
    Odrv4 I__4393 (
            .O(N__27665),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__4392 (
            .O(N__27658),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__4391 (
            .O(N__27653),
            .I(N__27650));
    InMux I__4390 (
            .O(N__27650),
            .I(N__27647));
    LocalMux I__4389 (
            .O(N__27647),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0 ));
    InMux I__4388 (
            .O(N__27644),
            .I(N__27641));
    LocalMux I__4387 (
            .O(N__27641),
            .I(\current_shift_inst.PI_CTRL.integrator_i_9 ));
    CascadeMux I__4386 (
            .O(N__27638),
            .I(N__27635));
    InMux I__4385 (
            .O(N__27635),
            .I(N__27631));
    InMux I__4384 (
            .O(N__27634),
            .I(N__27625));
    LocalMux I__4383 (
            .O(N__27631),
            .I(N__27622));
    InMux I__4382 (
            .O(N__27630),
            .I(N__27617));
    InMux I__4381 (
            .O(N__27629),
            .I(N__27617));
    InMux I__4380 (
            .O(N__27628),
            .I(N__27614));
    LocalMux I__4379 (
            .O(N__27625),
            .I(N__27611));
    Span4Mux_h I__4378 (
            .O(N__27622),
            .I(N__27608));
    LocalMux I__4377 (
            .O(N__27617),
            .I(N__27605));
    LocalMux I__4376 (
            .O(N__27614),
            .I(N__27602));
    Odrv4 I__4375 (
            .O(N__27611),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__4374 (
            .O(N__27608),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__4373 (
            .O(N__27605),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv12 I__4372 (
            .O(N__27602),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__4371 (
            .O(N__27593),
            .I(N__27590));
    InMux I__4370 (
            .O(N__27590),
            .I(N__27587));
    LocalMux I__4369 (
            .O(N__27587),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0 ));
    CascadeMux I__4368 (
            .O(N__27584),
            .I(N__27581));
    InMux I__4367 (
            .O(N__27581),
            .I(N__27578));
    LocalMux I__4366 (
            .O(N__27578),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0 ));
    InMux I__4365 (
            .O(N__27575),
            .I(N__27571));
    InMux I__4364 (
            .O(N__27574),
            .I(N__27568));
    LocalMux I__4363 (
            .O(N__27571),
            .I(N__27564));
    LocalMux I__4362 (
            .O(N__27568),
            .I(N__27561));
    InMux I__4361 (
            .O(N__27567),
            .I(N__27556));
    Span4Mux_h I__4360 (
            .O(N__27564),
            .I(N__27551));
    Span4Mux_h I__4359 (
            .O(N__27561),
            .I(N__27551));
    InMux I__4358 (
            .O(N__27560),
            .I(N__27546));
    InMux I__4357 (
            .O(N__27559),
            .I(N__27546));
    LocalMux I__4356 (
            .O(N__27556),
            .I(N__27543));
    Odrv4 I__4355 (
            .O(N__27551),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__4354 (
            .O(N__27546),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__4353 (
            .O(N__27543),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__4352 (
            .O(N__27536),
            .I(N__27533));
    LocalMux I__4351 (
            .O(N__27533),
            .I(\current_shift_inst.PI_CTRL.integrator_i_21 ));
    CascadeMux I__4350 (
            .O(N__27530),
            .I(N__27525));
    InMux I__4349 (
            .O(N__27529),
            .I(N__27522));
    InMux I__4348 (
            .O(N__27528),
            .I(N__27519));
    InMux I__4347 (
            .O(N__27525),
            .I(N__27515));
    LocalMux I__4346 (
            .O(N__27522),
            .I(N__27512));
    LocalMux I__4345 (
            .O(N__27519),
            .I(N__27509));
    InMux I__4344 (
            .O(N__27518),
            .I(N__27506));
    LocalMux I__4343 (
            .O(N__27515),
            .I(N__27503));
    Span4Mux_h I__4342 (
            .O(N__27512),
            .I(N__27500));
    Span4Mux_h I__4341 (
            .O(N__27509),
            .I(N__27496));
    LocalMux I__4340 (
            .O(N__27506),
            .I(N__27493));
    Span4Mux_v I__4339 (
            .O(N__27503),
            .I(N__27488));
    Span4Mux_v I__4338 (
            .O(N__27500),
            .I(N__27488));
    InMux I__4337 (
            .O(N__27499),
            .I(N__27485));
    Odrv4 I__4336 (
            .O(N__27496),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv12 I__4335 (
            .O(N__27493),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__4334 (
            .O(N__27488),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__4333 (
            .O(N__27485),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    CascadeMux I__4332 (
            .O(N__27476),
            .I(N__27473));
    InMux I__4331 (
            .O(N__27473),
            .I(N__27470));
    LocalMux I__4330 (
            .O(N__27470),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12 ));
    InMux I__4329 (
            .O(N__27467),
            .I(N__27464));
    LocalMux I__4328 (
            .O(N__27464),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0 ));
    CascadeMux I__4327 (
            .O(N__27461),
            .I(N__27458));
    InMux I__4326 (
            .O(N__27458),
            .I(N__27455));
    LocalMux I__4325 (
            .O(N__27455),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0 ));
    CascadeMux I__4324 (
            .O(N__27452),
            .I(N__27449));
    InMux I__4323 (
            .O(N__27449),
            .I(N__27446));
    LocalMux I__4322 (
            .O(N__27446),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0 ));
    CascadeMux I__4321 (
            .O(N__27443),
            .I(N__27440));
    InMux I__4320 (
            .O(N__27440),
            .I(N__27437));
    LocalMux I__4319 (
            .O(N__27437),
            .I(N__27434));
    Odrv4 I__4318 (
            .O(N__27434),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0 ));
    CascadeMux I__4317 (
            .O(N__27431),
            .I(N__27427));
    CascadeMux I__4316 (
            .O(N__27430),
            .I(N__27424));
    InMux I__4315 (
            .O(N__27427),
            .I(N__27419));
    InMux I__4314 (
            .O(N__27424),
            .I(N__27416));
    InMux I__4313 (
            .O(N__27423),
            .I(N__27413));
    InMux I__4312 (
            .O(N__27422),
            .I(N__27410));
    LocalMux I__4311 (
            .O(N__27419),
            .I(N__27404));
    LocalMux I__4310 (
            .O(N__27416),
            .I(N__27404));
    LocalMux I__4309 (
            .O(N__27413),
            .I(N__27401));
    LocalMux I__4308 (
            .O(N__27410),
            .I(N__27398));
    InMux I__4307 (
            .O(N__27409),
            .I(N__27395));
    Span4Mux_v I__4306 (
            .O(N__27404),
            .I(N__27388));
    Span4Mux_v I__4305 (
            .O(N__27401),
            .I(N__27388));
    Span4Mux_h I__4304 (
            .O(N__27398),
            .I(N__27388));
    LocalMux I__4303 (
            .O(N__27395),
            .I(N__27383));
    Span4Mux_h I__4302 (
            .O(N__27388),
            .I(N__27383));
    Odrv4 I__4301 (
            .O(N__27383),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__4300 (
            .O(N__27380),
            .I(N__27377));
    InMux I__4299 (
            .O(N__27377),
            .I(N__27374));
    LocalMux I__4298 (
            .O(N__27374),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0 ));
    InMux I__4297 (
            .O(N__27371),
            .I(N__27366));
    InMux I__4296 (
            .O(N__27370),
            .I(N__27362));
    CascadeMux I__4295 (
            .O(N__27369),
            .I(N__27359));
    LocalMux I__4294 (
            .O(N__27366),
            .I(N__27356));
    InMux I__4293 (
            .O(N__27365),
            .I(N__27353));
    LocalMux I__4292 (
            .O(N__27362),
            .I(N__27349));
    InMux I__4291 (
            .O(N__27359),
            .I(N__27346));
    Span4Mux_v I__4290 (
            .O(N__27356),
            .I(N__27341));
    LocalMux I__4289 (
            .O(N__27353),
            .I(N__27341));
    InMux I__4288 (
            .O(N__27352),
            .I(N__27338));
    Span4Mux_h I__4287 (
            .O(N__27349),
            .I(N__27335));
    LocalMux I__4286 (
            .O(N__27346),
            .I(N__27330));
    Span4Mux_h I__4285 (
            .O(N__27341),
            .I(N__27330));
    LocalMux I__4284 (
            .O(N__27338),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__4283 (
            .O(N__27335),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__4282 (
            .O(N__27330),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    CascadeMux I__4281 (
            .O(N__27323),
            .I(N__27320));
    InMux I__4280 (
            .O(N__27320),
            .I(N__27317));
    LocalMux I__4279 (
            .O(N__27317),
            .I(N__27314));
    Span4Mux_v I__4278 (
            .O(N__27314),
            .I(N__27311));
    Odrv4 I__4277 (
            .O(N__27311),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0 ));
    CascadeMux I__4276 (
            .O(N__27308),
            .I(N__27305));
    InMux I__4275 (
            .O(N__27305),
            .I(N__27302));
    LocalMux I__4274 (
            .O(N__27302),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0 ));
    InMux I__4273 (
            .O(N__27299),
            .I(N__27296));
    LocalMux I__4272 (
            .O(N__27296),
            .I(N__27293));
    Odrv4 I__4271 (
            .O(N__27293),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    CascadeMux I__4270 (
            .O(N__27290),
            .I(N__27287));
    InMux I__4269 (
            .O(N__27287),
            .I(N__27284));
    LocalMux I__4268 (
            .O(N__27284),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6 ));
    InMux I__4267 (
            .O(N__27281),
            .I(N__27278));
    LocalMux I__4266 (
            .O(N__27278),
            .I(\current_shift_inst.PI_CTRL.integrator_i_1 ));
    CascadeMux I__4265 (
            .O(N__27275),
            .I(N__27272));
    InMux I__4264 (
            .O(N__27272),
            .I(N__27268));
    InMux I__4263 (
            .O(N__27271),
            .I(N__27265));
    LocalMux I__4262 (
            .O(N__27268),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_14 ));
    LocalMux I__4261 (
            .O(N__27265),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_14 ));
    CascadeMux I__4260 (
            .O(N__27260),
            .I(N__27256));
    InMux I__4259 (
            .O(N__27259),
            .I(N__27253));
    InMux I__4258 (
            .O(N__27256),
            .I(N__27250));
    LocalMux I__4257 (
            .O(N__27253),
            .I(N__27247));
    LocalMux I__4256 (
            .O(N__27250),
            .I(N__27242));
    Span4Mux_h I__4255 (
            .O(N__27247),
            .I(N__27242));
    Span4Mux_h I__4254 (
            .O(N__27242),
            .I(N__27237));
    InMux I__4253 (
            .O(N__27241),
            .I(N__27232));
    InMux I__4252 (
            .O(N__27240),
            .I(N__27232));
    Odrv4 I__4251 (
            .O(N__27237),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__4250 (
            .O(N__27232),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__4249 (
            .O(N__27227),
            .I(N__27224));
    LocalMux I__4248 (
            .O(N__27224),
            .I(\current_shift_inst.PI_CTRL.integrator_i_2 ));
    CascadeMux I__4247 (
            .O(N__27221),
            .I(N__27218));
    InMux I__4246 (
            .O(N__27218),
            .I(N__27215));
    LocalMux I__4245 (
            .O(N__27215),
            .I(N__27212));
    Span4Mux_h I__4244 (
            .O(N__27212),
            .I(N__27209));
    Odrv4 I__4243 (
            .O(N__27209),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13 ));
    CascadeMux I__4242 (
            .O(N__27206),
            .I(N__27203));
    InMux I__4241 (
            .O(N__27203),
            .I(N__27197));
    InMux I__4240 (
            .O(N__27202),
            .I(N__27194));
    InMux I__4239 (
            .O(N__27201),
            .I(N__27190));
    InMux I__4238 (
            .O(N__27200),
            .I(N__27187));
    LocalMux I__4237 (
            .O(N__27197),
            .I(N__27184));
    LocalMux I__4236 (
            .O(N__27194),
            .I(N__27181));
    InMux I__4235 (
            .O(N__27193),
            .I(N__27178));
    LocalMux I__4234 (
            .O(N__27190),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__4233 (
            .O(N__27187),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv12 I__4232 (
            .O(N__27184),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__4231 (
            .O(N__27181),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__4230 (
            .O(N__27178),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__4229 (
            .O(N__27167),
            .I(N__27164));
    InMux I__4228 (
            .O(N__27164),
            .I(N__27161));
    LocalMux I__4227 (
            .O(N__27161),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8 ));
    CascadeMux I__4226 (
            .O(N__27158),
            .I(N__27154));
    InMux I__4225 (
            .O(N__27157),
            .I(N__27150));
    InMux I__4224 (
            .O(N__27154),
            .I(N__27146));
    InMux I__4223 (
            .O(N__27153),
            .I(N__27143));
    LocalMux I__4222 (
            .O(N__27150),
            .I(N__27140));
    InMux I__4221 (
            .O(N__27149),
            .I(N__27137));
    LocalMux I__4220 (
            .O(N__27146),
            .I(N__27132));
    LocalMux I__4219 (
            .O(N__27143),
            .I(N__27132));
    Span4Mux_h I__4218 (
            .O(N__27140),
            .I(N__27126));
    LocalMux I__4217 (
            .O(N__27137),
            .I(N__27126));
    Span4Mux_h I__4216 (
            .O(N__27132),
            .I(N__27123));
    InMux I__4215 (
            .O(N__27131),
            .I(N__27120));
    Odrv4 I__4214 (
            .O(N__27126),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__4213 (
            .O(N__27123),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__4212 (
            .O(N__27120),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    CascadeMux I__4211 (
            .O(N__27113),
            .I(N__27110));
    InMux I__4210 (
            .O(N__27110),
            .I(N__27107));
    LocalMux I__4209 (
            .O(N__27107),
            .I(\current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9 ));
    InMux I__4208 (
            .O(N__27104),
            .I(N__27100));
    CascadeMux I__4207 (
            .O(N__27103),
            .I(N__27097));
    LocalMux I__4206 (
            .O(N__27100),
            .I(N__27094));
    InMux I__4205 (
            .O(N__27097),
            .I(N__27091));
    Span4Mux_v I__4204 (
            .O(N__27094),
            .I(N__27088));
    LocalMux I__4203 (
            .O(N__27091),
            .I(N__27085));
    Span4Mux_h I__4202 (
            .O(N__27088),
            .I(N__27080));
    Span4Mux_v I__4201 (
            .O(N__27085),
            .I(N__27077));
    InMux I__4200 (
            .O(N__27084),
            .I(N__27072));
    InMux I__4199 (
            .O(N__27083),
            .I(N__27072));
    Odrv4 I__4198 (
            .O(N__27080),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__4197 (
            .O(N__27077),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__4196 (
            .O(N__27072),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__4195 (
            .O(N__27065),
            .I(N__27062));
    InMux I__4194 (
            .O(N__27062),
            .I(N__27059));
    LocalMux I__4193 (
            .O(N__27059),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5 ));
    CascadeMux I__4192 (
            .O(N__27056),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_ ));
    CascadeMux I__4191 (
            .O(N__27053),
            .I(N__27050));
    InMux I__4190 (
            .O(N__27050),
            .I(N__27045));
    InMux I__4189 (
            .O(N__27049),
            .I(N__27040));
    InMux I__4188 (
            .O(N__27048),
            .I(N__27040));
    LocalMux I__4187 (
            .O(N__27045),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__4186 (
            .O(N__27040),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__4185 (
            .O(N__27035),
            .I(N__27030));
    InMux I__4184 (
            .O(N__27034),
            .I(N__27025));
    InMux I__4183 (
            .O(N__27033),
            .I(N__27025));
    LocalMux I__4182 (
            .O(N__27030),
            .I(N__27022));
    LocalMux I__4181 (
            .O(N__27025),
            .I(N__27019));
    Span4Mux_h I__4180 (
            .O(N__27022),
            .I(N__27016));
    Span12Mux_h I__4179 (
            .O(N__27019),
            .I(N__27013));
    Span4Mux_v I__4178 (
            .O(N__27016),
            .I(N__27010));
    Span12Mux_v I__4177 (
            .O(N__27013),
            .I(N__27007));
    Span4Mux_v I__4176 (
            .O(N__27010),
            .I(N__27004));
    Odrv12 I__4175 (
            .O(N__27007),
            .I(il_min_comp2_c));
    Odrv4 I__4174 (
            .O(N__27004),
            .I(il_min_comp2_c));
    CascadeMux I__4173 (
            .O(N__26999),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2_cascade_ ));
    InMux I__4172 (
            .O(N__26996),
            .I(N__26993));
    LocalMux I__4171 (
            .O(N__26993),
            .I(N__26990));
    Sp12to4 I__4170 (
            .O(N__26990),
            .I(N__26984));
    InMux I__4169 (
            .O(N__26989),
            .I(N__26979));
    InMux I__4168 (
            .O(N__26988),
            .I(N__26979));
    InMux I__4167 (
            .O(N__26987),
            .I(N__26976));
    Odrv12 I__4166 (
            .O(N__26984),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__4165 (
            .O(N__26979),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__4164 (
            .O(N__26976),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__4163 (
            .O(N__26969),
            .I(N__26966));
    LocalMux I__4162 (
            .O(N__26966),
            .I(N__26963));
    Odrv4 I__4161 (
            .O(N__26963),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ));
    CascadeMux I__4160 (
            .O(N__26960),
            .I(N__26956));
    InMux I__4159 (
            .O(N__26959),
            .I(N__26953));
    InMux I__4158 (
            .O(N__26956),
            .I(N__26950));
    LocalMux I__4157 (
            .O(N__26953),
            .I(N__26945));
    LocalMux I__4156 (
            .O(N__26950),
            .I(N__26945));
    Span4Mux_h I__4155 (
            .O(N__26945),
            .I(N__26942));
    Span4Mux_h I__4154 (
            .O(N__26942),
            .I(N__26938));
    InMux I__4153 (
            .O(N__26941),
            .I(N__26935));
    Odrv4 I__4152 (
            .O(N__26938),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__4151 (
            .O(N__26935),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__4150 (
            .O(N__26930),
            .I(N__26927));
    LocalMux I__4149 (
            .O(N__26927),
            .I(N__26924));
    Odrv4 I__4148 (
            .O(N__26924),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    CascadeMux I__4147 (
            .O(N__26921),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0_cascade_ ));
    CascadeMux I__4146 (
            .O(N__26918),
            .I(N__26915));
    InMux I__4145 (
            .O(N__26915),
            .I(N__26912));
    LocalMux I__4144 (
            .O(N__26912),
            .I(N__26909));
    Span4Mux_v I__4143 (
            .O(N__26909),
            .I(N__26906));
    Odrv4 I__4142 (
            .O(N__26906),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4 ));
    InMux I__4141 (
            .O(N__26903),
            .I(N__26900));
    LocalMux I__4140 (
            .O(N__26900),
            .I(N__26897));
    Odrv4 I__4139 (
            .O(N__26897),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ));
    InMux I__4138 (
            .O(N__26894),
            .I(N__26891));
    LocalMux I__4137 (
            .O(N__26891),
            .I(N__26887));
    InMux I__4136 (
            .O(N__26890),
            .I(N__26884));
    Odrv12 I__4135 (
            .O(N__26887),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    LocalMux I__4134 (
            .O(N__26884),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    CascadeMux I__4133 (
            .O(N__26879),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_));
    InMux I__4132 (
            .O(N__26876),
            .I(N__26872));
    InMux I__4131 (
            .O(N__26875),
            .I(N__26869));
    LocalMux I__4130 (
            .O(N__26872),
            .I(N__26866));
    LocalMux I__4129 (
            .O(N__26869),
            .I(N__26861));
    Span4Mux_h I__4128 (
            .O(N__26866),
            .I(N__26858));
    InMux I__4127 (
            .O(N__26865),
            .I(N__26853));
    InMux I__4126 (
            .O(N__26864),
            .I(N__26853));
    Span4Mux_h I__4125 (
            .O(N__26861),
            .I(N__26850));
    Odrv4 I__4124 (
            .O(N__26858),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    LocalMux I__4123 (
            .O(N__26853),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__4122 (
            .O(N__26850),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    CascadeMux I__4121 (
            .O(N__26843),
            .I(N__26839));
    InMux I__4120 (
            .O(N__26842),
            .I(N__26834));
    InMux I__4119 (
            .O(N__26839),
            .I(N__26834));
    LocalMux I__4118 (
            .O(N__26834),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ));
    InMux I__4117 (
            .O(N__26831),
            .I(N__26828));
    LocalMux I__4116 (
            .O(N__26828),
            .I(N__26823));
    InMux I__4115 (
            .O(N__26827),
            .I(N__26820));
    InMux I__4114 (
            .O(N__26826),
            .I(N__26817));
    Span4Mux_v I__4113 (
            .O(N__26823),
            .I(N__26814));
    LocalMux I__4112 (
            .O(N__26820),
            .I(N__26811));
    LocalMux I__4111 (
            .O(N__26817),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv4 I__4110 (
            .O(N__26814),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv12 I__4109 (
            .O(N__26811),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    InMux I__4108 (
            .O(N__26804),
            .I(N__26798));
    InMux I__4107 (
            .O(N__26803),
            .I(N__26798));
    LocalMux I__4106 (
            .O(N__26798),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ));
    InMux I__4105 (
            .O(N__26795),
            .I(N__26792));
    LocalMux I__4104 (
            .O(N__26792),
            .I(N__26788));
    InMux I__4103 (
            .O(N__26791),
            .I(N__26782));
    Span4Mux_h I__4102 (
            .O(N__26788),
            .I(N__26779));
    InMux I__4101 (
            .O(N__26787),
            .I(N__26772));
    InMux I__4100 (
            .O(N__26786),
            .I(N__26772));
    InMux I__4099 (
            .O(N__26785),
            .I(N__26772));
    LocalMux I__4098 (
            .O(N__26782),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__4097 (
            .O(N__26779),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__4096 (
            .O(N__26772),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    CascadeMux I__4095 (
            .O(N__26765),
            .I(N__26762));
    InMux I__4094 (
            .O(N__26762),
            .I(N__26759));
    LocalMux I__4093 (
            .O(N__26759),
            .I(N__26755));
    InMux I__4092 (
            .O(N__26758),
            .I(N__26752));
    Span4Mux_v I__4091 (
            .O(N__26755),
            .I(N__26749));
    LocalMux I__4090 (
            .O(N__26752),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__4089 (
            .O(N__26749),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    CascadeMux I__4088 (
            .O(N__26744),
            .I(N__26740));
    InMux I__4087 (
            .O(N__26743),
            .I(N__26737));
    InMux I__4086 (
            .O(N__26740),
            .I(N__26733));
    LocalMux I__4085 (
            .O(N__26737),
            .I(N__26730));
    InMux I__4084 (
            .O(N__26736),
            .I(N__26725));
    LocalMux I__4083 (
            .O(N__26733),
            .I(N__26722));
    Span4Mux_h I__4082 (
            .O(N__26730),
            .I(N__26719));
    InMux I__4081 (
            .O(N__26729),
            .I(N__26714));
    InMux I__4080 (
            .O(N__26728),
            .I(N__26714));
    LocalMux I__4079 (
            .O(N__26725),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    Odrv4 I__4078 (
            .O(N__26722),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    Odrv4 I__4077 (
            .O(N__26719),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__4076 (
            .O(N__26714),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__4075 (
            .O(N__26705),
            .I(N__26696));
    InMux I__4074 (
            .O(N__26704),
            .I(N__26696));
    InMux I__4073 (
            .O(N__26703),
            .I(N__26696));
    LocalMux I__4072 (
            .O(N__26696),
            .I(\phase_controller_inst2.tr_time_passed ));
    CascadeMux I__4071 (
            .O(N__26693),
            .I(N__26690));
    InMux I__4070 (
            .O(N__26690),
            .I(N__26686));
    InMux I__4069 (
            .O(N__26689),
            .I(N__26683));
    LocalMux I__4068 (
            .O(N__26686),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__4067 (
            .O(N__26683),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__4066 (
            .O(N__26678),
            .I(N__26675));
    LocalMux I__4065 (
            .O(N__26675),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    InMux I__4064 (
            .O(N__26672),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__4063 (
            .O(N__26669),
            .I(N__26666));
    InMux I__4062 (
            .O(N__26666),
            .I(N__26662));
    InMux I__4061 (
            .O(N__26665),
            .I(N__26659));
    LocalMux I__4060 (
            .O(N__26662),
            .I(N__26653));
    LocalMux I__4059 (
            .O(N__26659),
            .I(N__26653));
    InMux I__4058 (
            .O(N__26658),
            .I(N__26650));
    Span4Mux_v I__4057 (
            .O(N__26653),
            .I(N__26647));
    LocalMux I__4056 (
            .O(N__26650),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__4055 (
            .O(N__26647),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__4054 (
            .O(N__26642),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__4053 (
            .O(N__26639),
            .I(N__26635));
    CascadeMux I__4052 (
            .O(N__26638),
            .I(N__26632));
    InMux I__4051 (
            .O(N__26635),
            .I(N__26629));
    InMux I__4050 (
            .O(N__26632),
            .I(N__26626));
    LocalMux I__4049 (
            .O(N__26629),
            .I(N__26620));
    LocalMux I__4048 (
            .O(N__26626),
            .I(N__26620));
    InMux I__4047 (
            .O(N__26625),
            .I(N__26617));
    Span4Mux_v I__4046 (
            .O(N__26620),
            .I(N__26614));
    LocalMux I__4045 (
            .O(N__26617),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__4044 (
            .O(N__26614),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__4043 (
            .O(N__26609),
            .I(bfn_9_11_0_));
    CascadeMux I__4042 (
            .O(N__26606),
            .I(N__26603));
    InMux I__4041 (
            .O(N__26603),
            .I(N__26598));
    InMux I__4040 (
            .O(N__26602),
            .I(N__26595));
    InMux I__4039 (
            .O(N__26601),
            .I(N__26592));
    LocalMux I__4038 (
            .O(N__26598),
            .I(N__26587));
    LocalMux I__4037 (
            .O(N__26595),
            .I(N__26587));
    LocalMux I__4036 (
            .O(N__26592),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv12 I__4035 (
            .O(N__26587),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__4034 (
            .O(N__26582),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__4033 (
            .O(N__26579),
            .I(N__26572));
    InMux I__4032 (
            .O(N__26578),
            .I(N__26572));
    InMux I__4031 (
            .O(N__26577),
            .I(N__26569));
    LocalMux I__4030 (
            .O(N__26572),
            .I(N__26566));
    LocalMux I__4029 (
            .O(N__26569),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv12 I__4028 (
            .O(N__26566),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    CascadeMux I__4027 (
            .O(N__26561),
            .I(N__26558));
    InMux I__4026 (
            .O(N__26558),
            .I(N__26554));
    InMux I__4025 (
            .O(N__26557),
            .I(N__26551));
    LocalMux I__4024 (
            .O(N__26554),
            .I(N__26548));
    LocalMux I__4023 (
            .O(N__26551),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv12 I__4022 (
            .O(N__26548),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__4021 (
            .O(N__26543),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__4020 (
            .O(N__26540),
            .I(N__26537));
    LocalMux I__4019 (
            .O(N__26537),
            .I(N__26533));
    InMux I__4018 (
            .O(N__26536),
            .I(N__26530));
    Span4Mux_v I__4017 (
            .O(N__26533),
            .I(N__26527));
    LocalMux I__4016 (
            .O(N__26530),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__4015 (
            .O(N__26527),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__4014 (
            .O(N__26522),
            .I(N__26519));
    InMux I__4013 (
            .O(N__26519),
            .I(N__26514));
    InMux I__4012 (
            .O(N__26518),
            .I(N__26511));
    InMux I__4011 (
            .O(N__26517),
            .I(N__26508));
    LocalMux I__4010 (
            .O(N__26514),
            .I(N__26503));
    LocalMux I__4009 (
            .O(N__26511),
            .I(N__26503));
    LocalMux I__4008 (
            .O(N__26508),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv12 I__4007 (
            .O(N__26503),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__4006 (
            .O(N__26498),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__4005 (
            .O(N__26495),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__4004 (
            .O(N__26492),
            .I(N__26487));
    CEMux I__4003 (
            .O(N__26491),
            .I(N__26484));
    CEMux I__4002 (
            .O(N__26490),
            .I(N__26480));
    LocalMux I__4001 (
            .O(N__26487),
            .I(N__26476));
    LocalMux I__4000 (
            .O(N__26484),
            .I(N__26473));
    CEMux I__3999 (
            .O(N__26483),
            .I(N__26470));
    LocalMux I__3998 (
            .O(N__26480),
            .I(N__26467));
    CEMux I__3997 (
            .O(N__26479),
            .I(N__26464));
    Span4Mux_v I__3996 (
            .O(N__26476),
            .I(N__26457));
    Span4Mux_v I__3995 (
            .O(N__26473),
            .I(N__26457));
    LocalMux I__3994 (
            .O(N__26470),
            .I(N__26457));
    Span4Mux_h I__3993 (
            .O(N__26467),
            .I(N__26454));
    LocalMux I__3992 (
            .O(N__26464),
            .I(N__26451));
    Odrv4 I__3991 (
            .O(N__26457),
            .I(\delay_measurement_inst.delay_tr_timer.N_203_i ));
    Odrv4 I__3990 (
            .O(N__26454),
            .I(\delay_measurement_inst.delay_tr_timer.N_203_i ));
    Odrv4 I__3989 (
            .O(N__26451),
            .I(\delay_measurement_inst.delay_tr_timer.N_203_i ));
    InMux I__3988 (
            .O(N__26444),
            .I(N__26440));
    InMux I__3987 (
            .O(N__26443),
            .I(N__26437));
    LocalMux I__3986 (
            .O(N__26440),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    LocalMux I__3985 (
            .O(N__26437),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    InMux I__3984 (
            .O(N__26432),
            .I(N__26428));
    InMux I__3983 (
            .O(N__26431),
            .I(N__26425));
    LocalMux I__3982 (
            .O(N__26428),
            .I(N__26420));
    LocalMux I__3981 (
            .O(N__26425),
            .I(N__26417));
    InMux I__3980 (
            .O(N__26424),
            .I(N__26412));
    InMux I__3979 (
            .O(N__26423),
            .I(N__26412));
    Span4Mux_v I__3978 (
            .O(N__26420),
            .I(N__26407));
    Span4Mux_h I__3977 (
            .O(N__26417),
            .I(N__26407));
    LocalMux I__3976 (
            .O(N__26412),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__3975 (
            .O(N__26407),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    CascadeMux I__3974 (
            .O(N__26402),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_));
    InMux I__3973 (
            .O(N__26399),
            .I(N__26393));
    InMux I__3972 (
            .O(N__26398),
            .I(N__26393));
    LocalMux I__3971 (
            .O(N__26393),
            .I(N__26389));
    InMux I__3970 (
            .O(N__26392),
            .I(N__26386));
    Span4Mux_v I__3969 (
            .O(N__26389),
            .I(N__26383));
    LocalMux I__3968 (
            .O(N__26386),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__3967 (
            .O(N__26383),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__3966 (
            .O(N__26378),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__3965 (
            .O(N__26375),
            .I(N__26371));
    CascadeMux I__3964 (
            .O(N__26374),
            .I(N__26368));
    InMux I__3963 (
            .O(N__26371),
            .I(N__26362));
    InMux I__3962 (
            .O(N__26368),
            .I(N__26362));
    InMux I__3961 (
            .O(N__26367),
            .I(N__26359));
    LocalMux I__3960 (
            .O(N__26362),
            .I(N__26356));
    LocalMux I__3959 (
            .O(N__26359),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv12 I__3958 (
            .O(N__26356),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__3957 (
            .O(N__26351),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__3956 (
            .O(N__26348),
            .I(N__26344));
    CascadeMux I__3955 (
            .O(N__26347),
            .I(N__26341));
    InMux I__3954 (
            .O(N__26344),
            .I(N__26338));
    InMux I__3953 (
            .O(N__26341),
            .I(N__26335));
    LocalMux I__3952 (
            .O(N__26338),
            .I(N__26329));
    LocalMux I__3951 (
            .O(N__26335),
            .I(N__26329));
    InMux I__3950 (
            .O(N__26334),
            .I(N__26326));
    Span4Mux_v I__3949 (
            .O(N__26329),
            .I(N__26323));
    LocalMux I__3948 (
            .O(N__26326),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__3947 (
            .O(N__26323),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__3946 (
            .O(N__26318),
            .I(bfn_9_10_0_));
    CascadeMux I__3945 (
            .O(N__26315),
            .I(N__26312));
    InMux I__3944 (
            .O(N__26312),
            .I(N__26309));
    LocalMux I__3943 (
            .O(N__26309),
            .I(N__26304));
    InMux I__3942 (
            .O(N__26308),
            .I(N__26301));
    InMux I__3941 (
            .O(N__26307),
            .I(N__26298));
    Sp12to4 I__3940 (
            .O(N__26304),
            .I(N__26293));
    LocalMux I__3939 (
            .O(N__26301),
            .I(N__26293));
    LocalMux I__3938 (
            .O(N__26298),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv12 I__3937 (
            .O(N__26293),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__3936 (
            .O(N__26288),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__3935 (
            .O(N__26285),
            .I(N__26278));
    InMux I__3934 (
            .O(N__26284),
            .I(N__26278));
    InMux I__3933 (
            .O(N__26283),
            .I(N__26275));
    LocalMux I__3932 (
            .O(N__26278),
            .I(N__26272));
    LocalMux I__3931 (
            .O(N__26275),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv12 I__3930 (
            .O(N__26272),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__3929 (
            .O(N__26267),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__3928 (
            .O(N__26264),
            .I(N__26257));
    InMux I__3927 (
            .O(N__26263),
            .I(N__26257));
    InMux I__3926 (
            .O(N__26262),
            .I(N__26254));
    LocalMux I__3925 (
            .O(N__26257),
            .I(N__26251));
    LocalMux I__3924 (
            .O(N__26254),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv12 I__3923 (
            .O(N__26251),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__3922 (
            .O(N__26246),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__3921 (
            .O(N__26243),
            .I(N__26239));
    CascadeMux I__3920 (
            .O(N__26242),
            .I(N__26236));
    InMux I__3919 (
            .O(N__26239),
            .I(N__26230));
    InMux I__3918 (
            .O(N__26236),
            .I(N__26230));
    InMux I__3917 (
            .O(N__26235),
            .I(N__26227));
    LocalMux I__3916 (
            .O(N__26230),
            .I(N__26224));
    LocalMux I__3915 (
            .O(N__26227),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv12 I__3914 (
            .O(N__26224),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__3913 (
            .O(N__26219),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__3912 (
            .O(N__26216),
            .I(N__26212));
    CascadeMux I__3911 (
            .O(N__26215),
            .I(N__26209));
    InMux I__3910 (
            .O(N__26212),
            .I(N__26203));
    InMux I__3909 (
            .O(N__26209),
            .I(N__26203));
    InMux I__3908 (
            .O(N__26208),
            .I(N__26200));
    LocalMux I__3907 (
            .O(N__26203),
            .I(N__26197));
    LocalMux I__3906 (
            .O(N__26200),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv12 I__3905 (
            .O(N__26197),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__3904 (
            .O(N__26192),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__3903 (
            .O(N__26189),
            .I(N__26183));
    InMux I__3902 (
            .O(N__26188),
            .I(N__26183));
    LocalMux I__3901 (
            .O(N__26183),
            .I(N__26179));
    InMux I__3900 (
            .O(N__26182),
            .I(N__26176));
    Span4Mux_v I__3899 (
            .O(N__26179),
            .I(N__26173));
    LocalMux I__3898 (
            .O(N__26176),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__3897 (
            .O(N__26173),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__3896 (
            .O(N__26168),
            .I(N__26162));
    InMux I__3895 (
            .O(N__26167),
            .I(N__26162));
    LocalMux I__3894 (
            .O(N__26162),
            .I(N__26158));
    InMux I__3893 (
            .O(N__26161),
            .I(N__26155));
    Span4Mux_v I__3892 (
            .O(N__26158),
            .I(N__26152));
    LocalMux I__3891 (
            .O(N__26155),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__3890 (
            .O(N__26152),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__3889 (
            .O(N__26147),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__3888 (
            .O(N__26144),
            .I(N__26138));
    InMux I__3887 (
            .O(N__26143),
            .I(N__26138));
    LocalMux I__3886 (
            .O(N__26138),
            .I(N__26134));
    InMux I__3885 (
            .O(N__26137),
            .I(N__26131));
    Span4Mux_v I__3884 (
            .O(N__26134),
            .I(N__26128));
    LocalMux I__3883 (
            .O(N__26131),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__3882 (
            .O(N__26128),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__3881 (
            .O(N__26123),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__3880 (
            .O(N__26120),
            .I(N__26116));
    CascadeMux I__3879 (
            .O(N__26119),
            .I(N__26113));
    InMux I__3878 (
            .O(N__26116),
            .I(N__26110));
    InMux I__3877 (
            .O(N__26113),
            .I(N__26107));
    LocalMux I__3876 (
            .O(N__26110),
            .I(N__26101));
    LocalMux I__3875 (
            .O(N__26107),
            .I(N__26101));
    InMux I__3874 (
            .O(N__26106),
            .I(N__26098));
    Span4Mux_v I__3873 (
            .O(N__26101),
            .I(N__26095));
    LocalMux I__3872 (
            .O(N__26098),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__3871 (
            .O(N__26095),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__3870 (
            .O(N__26090),
            .I(bfn_9_9_0_));
    CascadeMux I__3869 (
            .O(N__26087),
            .I(N__26083));
    CascadeMux I__3868 (
            .O(N__26086),
            .I(N__26080));
    InMux I__3867 (
            .O(N__26083),
            .I(N__26076));
    InMux I__3866 (
            .O(N__26080),
            .I(N__26073));
    InMux I__3865 (
            .O(N__26079),
            .I(N__26070));
    LocalMux I__3864 (
            .O(N__26076),
            .I(N__26065));
    LocalMux I__3863 (
            .O(N__26073),
            .I(N__26065));
    LocalMux I__3862 (
            .O(N__26070),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv12 I__3861 (
            .O(N__26065),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__3860 (
            .O(N__26060),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__3859 (
            .O(N__26057),
            .I(N__26051));
    InMux I__3858 (
            .O(N__26056),
            .I(N__26051));
    LocalMux I__3857 (
            .O(N__26051),
            .I(N__26047));
    InMux I__3856 (
            .O(N__26050),
            .I(N__26044));
    Span4Mux_v I__3855 (
            .O(N__26047),
            .I(N__26041));
    LocalMux I__3854 (
            .O(N__26044),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__3853 (
            .O(N__26041),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__3852 (
            .O(N__26036),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__3851 (
            .O(N__26033),
            .I(N__26030));
    InMux I__3850 (
            .O(N__26030),
            .I(N__26026));
    InMux I__3849 (
            .O(N__26029),
            .I(N__26023));
    LocalMux I__3848 (
            .O(N__26026),
            .I(N__26017));
    LocalMux I__3847 (
            .O(N__26023),
            .I(N__26017));
    InMux I__3846 (
            .O(N__26022),
            .I(N__26014));
    Span4Mux_v I__3845 (
            .O(N__26017),
            .I(N__26011));
    LocalMux I__3844 (
            .O(N__26014),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__3843 (
            .O(N__26011),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__3842 (
            .O(N__26006),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__3841 (
            .O(N__26003),
            .I(N__25999));
    CascadeMux I__3840 (
            .O(N__26002),
            .I(N__25996));
    InMux I__3839 (
            .O(N__25999),
            .I(N__25990));
    InMux I__3838 (
            .O(N__25996),
            .I(N__25990));
    InMux I__3837 (
            .O(N__25995),
            .I(N__25987));
    LocalMux I__3836 (
            .O(N__25990),
            .I(N__25984));
    LocalMux I__3835 (
            .O(N__25987),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv12 I__3834 (
            .O(N__25984),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__3833 (
            .O(N__25979),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__3832 (
            .O(N__25976),
            .I(N__25969));
    InMux I__3831 (
            .O(N__25975),
            .I(N__25969));
    InMux I__3830 (
            .O(N__25974),
            .I(N__25966));
    LocalMux I__3829 (
            .O(N__25969),
            .I(N__25963));
    LocalMux I__3828 (
            .O(N__25966),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv12 I__3827 (
            .O(N__25963),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__3826 (
            .O(N__25958),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__3825 (
            .O(N__25955),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__3824 (
            .O(N__25952),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__3823 (
            .O(N__25949),
            .I(N__25911));
    InMux I__3822 (
            .O(N__25948),
            .I(N__25911));
    InMux I__3821 (
            .O(N__25947),
            .I(N__25911));
    InMux I__3820 (
            .O(N__25946),
            .I(N__25911));
    InMux I__3819 (
            .O(N__25945),
            .I(N__25902));
    InMux I__3818 (
            .O(N__25944),
            .I(N__25902));
    InMux I__3817 (
            .O(N__25943),
            .I(N__25902));
    InMux I__3816 (
            .O(N__25942),
            .I(N__25902));
    InMux I__3815 (
            .O(N__25941),
            .I(N__25893));
    InMux I__3814 (
            .O(N__25940),
            .I(N__25893));
    InMux I__3813 (
            .O(N__25939),
            .I(N__25893));
    InMux I__3812 (
            .O(N__25938),
            .I(N__25893));
    InMux I__3811 (
            .O(N__25937),
            .I(N__25888));
    InMux I__3810 (
            .O(N__25936),
            .I(N__25888));
    InMux I__3809 (
            .O(N__25935),
            .I(N__25879));
    InMux I__3808 (
            .O(N__25934),
            .I(N__25879));
    InMux I__3807 (
            .O(N__25933),
            .I(N__25879));
    InMux I__3806 (
            .O(N__25932),
            .I(N__25879));
    InMux I__3805 (
            .O(N__25931),
            .I(N__25870));
    InMux I__3804 (
            .O(N__25930),
            .I(N__25870));
    InMux I__3803 (
            .O(N__25929),
            .I(N__25870));
    InMux I__3802 (
            .O(N__25928),
            .I(N__25870));
    InMux I__3801 (
            .O(N__25927),
            .I(N__25861));
    InMux I__3800 (
            .O(N__25926),
            .I(N__25861));
    InMux I__3799 (
            .O(N__25925),
            .I(N__25861));
    InMux I__3798 (
            .O(N__25924),
            .I(N__25861));
    InMux I__3797 (
            .O(N__25923),
            .I(N__25852));
    InMux I__3796 (
            .O(N__25922),
            .I(N__25852));
    InMux I__3795 (
            .O(N__25921),
            .I(N__25852));
    InMux I__3794 (
            .O(N__25920),
            .I(N__25852));
    LocalMux I__3793 (
            .O(N__25911),
            .I(N__25845));
    LocalMux I__3792 (
            .O(N__25902),
            .I(N__25845));
    LocalMux I__3791 (
            .O(N__25893),
            .I(N__25845));
    LocalMux I__3790 (
            .O(N__25888),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__3789 (
            .O(N__25879),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__3788 (
            .O(N__25870),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__3787 (
            .O(N__25861),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__3786 (
            .O(N__25852),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__3785 (
            .O(N__25845),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__3784 (
            .O(N__25832),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__3783 (
            .O(N__25829),
            .I(N__25826));
    LocalMux I__3782 (
            .O(N__25826),
            .I(N__25822));
    CEMux I__3781 (
            .O(N__25825),
            .I(N__25819));
    Span4Mux_v I__3780 (
            .O(N__25822),
            .I(N__25813));
    LocalMux I__3779 (
            .O(N__25819),
            .I(N__25813));
    CEMux I__3778 (
            .O(N__25818),
            .I(N__25810));
    Span4Mux_v I__3777 (
            .O(N__25813),
            .I(N__25806));
    LocalMux I__3776 (
            .O(N__25810),
            .I(N__25803));
    CEMux I__3775 (
            .O(N__25809),
            .I(N__25800));
    Span4Mux_h I__3774 (
            .O(N__25806),
            .I(N__25795));
    Span4Mux_v I__3773 (
            .O(N__25803),
            .I(N__25795));
    LocalMux I__3772 (
            .O(N__25800),
            .I(N__25792));
    Odrv4 I__3771 (
            .O(N__25795),
            .I(\delay_measurement_inst.delay_tr_timer.N_204_i ));
    Odrv12 I__3770 (
            .O(N__25792),
            .I(\delay_measurement_inst.delay_tr_timer.N_204_i ));
    CascadeMux I__3769 (
            .O(N__25787),
            .I(N__25783));
    InMux I__3768 (
            .O(N__25786),
            .I(N__25780));
    InMux I__3767 (
            .O(N__25783),
            .I(N__25777));
    LocalMux I__3766 (
            .O(N__25780),
            .I(N__25771));
    LocalMux I__3765 (
            .O(N__25777),
            .I(N__25771));
    InMux I__3764 (
            .O(N__25776),
            .I(N__25768));
    Span4Mux_v I__3763 (
            .O(N__25771),
            .I(N__25765));
    LocalMux I__3762 (
            .O(N__25768),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__3761 (
            .O(N__25765),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__3760 (
            .O(N__25760),
            .I(N__25757));
    LocalMux I__3759 (
            .O(N__25757),
            .I(N__25753));
    InMux I__3758 (
            .O(N__25756),
            .I(N__25750));
    Sp12to4 I__3757 (
            .O(N__25753),
            .I(N__25744));
    LocalMux I__3756 (
            .O(N__25750),
            .I(N__25744));
    InMux I__3755 (
            .O(N__25749),
            .I(N__25741));
    Odrv12 I__3754 (
            .O(N__25744),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__3753 (
            .O(N__25741),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__3752 (
            .O(N__25736),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__3751 (
            .O(N__25733),
            .I(N__25727));
    InMux I__3750 (
            .O(N__25732),
            .I(N__25727));
    LocalMux I__3749 (
            .O(N__25727),
            .I(N__25723));
    InMux I__3748 (
            .O(N__25726),
            .I(N__25720));
    Span4Mux_v I__3747 (
            .O(N__25723),
            .I(N__25717));
    LocalMux I__3746 (
            .O(N__25720),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__3745 (
            .O(N__25717),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__3744 (
            .O(N__25712),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__3743 (
            .O(N__25709),
            .I(N__25705));
    InMux I__3742 (
            .O(N__25708),
            .I(N__25702));
    InMux I__3741 (
            .O(N__25705),
            .I(N__25699));
    LocalMux I__3740 (
            .O(N__25702),
            .I(N__25695));
    LocalMux I__3739 (
            .O(N__25699),
            .I(N__25692));
    InMux I__3738 (
            .O(N__25698),
            .I(N__25689));
    Span4Mux_v I__3737 (
            .O(N__25695),
            .I(N__25684));
    Span4Mux_v I__3736 (
            .O(N__25692),
            .I(N__25684));
    LocalMux I__3735 (
            .O(N__25689),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__3734 (
            .O(N__25684),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__3733 (
            .O(N__25679),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__3732 (
            .O(N__25676),
            .I(N__25672));
    CascadeMux I__3731 (
            .O(N__25675),
            .I(N__25669));
    InMux I__3730 (
            .O(N__25672),
            .I(N__25663));
    InMux I__3729 (
            .O(N__25669),
            .I(N__25663));
    InMux I__3728 (
            .O(N__25668),
            .I(N__25660));
    LocalMux I__3727 (
            .O(N__25663),
            .I(N__25657));
    LocalMux I__3726 (
            .O(N__25660),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv12 I__3725 (
            .O(N__25657),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__3724 (
            .O(N__25652),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__3723 (
            .O(N__25649),
            .I(N__25645));
    CascadeMux I__3722 (
            .O(N__25648),
            .I(N__25642));
    InMux I__3721 (
            .O(N__25645),
            .I(N__25636));
    InMux I__3720 (
            .O(N__25642),
            .I(N__25636));
    InMux I__3719 (
            .O(N__25641),
            .I(N__25633));
    LocalMux I__3718 (
            .O(N__25636),
            .I(N__25630));
    LocalMux I__3717 (
            .O(N__25633),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv12 I__3716 (
            .O(N__25630),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__3715 (
            .O(N__25625),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__3714 (
            .O(N__25622),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__3713 (
            .O(N__25619),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__3712 (
            .O(N__25616),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__3711 (
            .O(N__25613),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__3710 (
            .O(N__25610),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__3709 (
            .O(N__25607),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__3708 (
            .O(N__25604),
            .I(bfn_9_7_0_));
    InMux I__3707 (
            .O(N__25601),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__3706 (
            .O(N__25598),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__3705 (
            .O(N__25595),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__3704 (
            .O(N__25592),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__3703 (
            .O(N__25589),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__3702 (
            .O(N__25586),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__3701 (
            .O(N__25583),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__3700 (
            .O(N__25580),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__3699 (
            .O(N__25577),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__3698 (
            .O(N__25574),
            .I(bfn_9_6_0_));
    InMux I__3697 (
            .O(N__25571),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__3696 (
            .O(N__25568),
            .I(bfn_9_4_0_));
    InMux I__3695 (
            .O(N__25565),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__3694 (
            .O(N__25562),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__3693 (
            .O(N__25559),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__3692 (
            .O(N__25556),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__3691 (
            .O(N__25553),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__3690 (
            .O(N__25550),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__3689 (
            .O(N__25547),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__3688 (
            .O(N__25544),
            .I(bfn_9_5_0_));
    InMux I__3687 (
            .O(N__25541),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ));
    InMux I__3686 (
            .O(N__25538),
            .I(N__25535));
    LocalMux I__3685 (
            .O(N__25535),
            .I(N__25532));
    Odrv4 I__3684 (
            .O(N__25532),
            .I(\current_shift_inst.PI_CTRL.integrator_i_30 ));
    InMux I__3683 (
            .O(N__25529),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ));
    InMux I__3682 (
            .O(N__25526),
            .I(bfn_8_20_0_));
    InMux I__3681 (
            .O(N__25523),
            .I(N__25520));
    LocalMux I__3680 (
            .O(N__25520),
            .I(\current_shift_inst.PI_CTRL.integrator_i_24 ));
    InMux I__3679 (
            .O(N__25517),
            .I(N__25514));
    LocalMux I__3678 (
            .O(N__25514),
            .I(\current_shift_inst.PI_CTRL.integrator_i_26 ));
    InMux I__3677 (
            .O(N__25511),
            .I(N__25508));
    LocalMux I__3676 (
            .O(N__25508),
            .I(N__25505));
    Odrv4 I__3675 (
            .O(N__25505),
            .I(\current_shift_inst.PI_CTRL.integrator_i_25 ));
    CascadeMux I__3674 (
            .O(N__25502),
            .I(N__25499));
    InMux I__3673 (
            .O(N__25499),
            .I(N__25495));
    InMux I__3672 (
            .O(N__25498),
            .I(N__25492));
    LocalMux I__3671 (
            .O(N__25495),
            .I(N__25488));
    LocalMux I__3670 (
            .O(N__25492),
            .I(N__25484));
    InMux I__3669 (
            .O(N__25491),
            .I(N__25481));
    Span4Mux_v I__3668 (
            .O(N__25488),
            .I(N__25478));
    InMux I__3667 (
            .O(N__25487),
            .I(N__25475));
    Span4Mux_v I__3666 (
            .O(N__25484),
            .I(N__25472));
    LocalMux I__3665 (
            .O(N__25481),
            .I(N__25469));
    Odrv4 I__3664 (
            .O(N__25478),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__3663 (
            .O(N__25475),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__3662 (
            .O(N__25472),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__3661 (
            .O(N__25469),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__3660 (
            .O(N__25460),
            .I(N__25457));
    LocalMux I__3659 (
            .O(N__25457),
            .I(\current_shift_inst.PI_CTRL.integrator_i_28 ));
    InMux I__3658 (
            .O(N__25454),
            .I(N__25451));
    LocalMux I__3657 (
            .O(N__25451),
            .I(N__25448));
    Odrv4 I__3656 (
            .O(N__25448),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    IoInMux I__3655 (
            .O(N__25445),
            .I(N__25442));
    LocalMux I__3654 (
            .O(N__25442),
            .I(N__25439));
    Odrv12 I__3653 (
            .O(N__25439),
            .I(s4_phy_c));
    CascadeMux I__3652 (
            .O(N__25436),
            .I(N__25433));
    InMux I__3651 (
            .O(N__25433),
            .I(N__25430));
    LocalMux I__3650 (
            .O(N__25430),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__3649 (
            .O(N__25427),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ));
    InMux I__3648 (
            .O(N__25424),
            .I(N__25421));
    LocalMux I__3647 (
            .O(N__25421),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__3646 (
            .O(N__25418),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ));
    CascadeMux I__3645 (
            .O(N__25415),
            .I(N__25412));
    InMux I__3644 (
            .O(N__25412),
            .I(N__25409));
    LocalMux I__3643 (
            .O(N__25409),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__3642 (
            .O(N__25406),
            .I(bfn_8_19_0_));
    InMux I__3641 (
            .O(N__25403),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ));
    CascadeMux I__3640 (
            .O(N__25400),
            .I(N__25397));
    InMux I__3639 (
            .O(N__25397),
            .I(N__25394));
    LocalMux I__3638 (
            .O(N__25394),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__3637 (
            .O(N__25391),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ));
    CascadeMux I__3636 (
            .O(N__25388),
            .I(N__25385));
    InMux I__3635 (
            .O(N__25385),
            .I(N__25382));
    LocalMux I__3634 (
            .O(N__25382),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__3633 (
            .O(N__25379),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ));
    InMux I__3632 (
            .O(N__25376),
            .I(N__25373));
    LocalMux I__3631 (
            .O(N__25373),
            .I(N__25370));
    Odrv4 I__3630 (
            .O(N__25370),
            .I(\current_shift_inst.PI_CTRL.integrator_i_27 ));
    InMux I__3629 (
            .O(N__25367),
            .I(N__25364));
    LocalMux I__3628 (
            .O(N__25364),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__3627 (
            .O(N__25361),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ));
    InMux I__3626 (
            .O(N__25358),
            .I(N__25355));
    LocalMux I__3625 (
            .O(N__25355),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__3624 (
            .O(N__25352),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ));
    InMux I__3623 (
            .O(N__25349),
            .I(N__25346));
    LocalMux I__3622 (
            .O(N__25346),
            .I(N__25343));
    Odrv12 I__3621 (
            .O(N__25343),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__3620 (
            .O(N__25340),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ));
    InMux I__3619 (
            .O(N__25337),
            .I(N__25334));
    LocalMux I__3618 (
            .O(N__25334),
            .I(N__25331));
    Odrv12 I__3617 (
            .O(N__25331),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__3616 (
            .O(N__25328),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ));
    InMux I__3615 (
            .O(N__25325),
            .I(N__25322));
    LocalMux I__3614 (
            .O(N__25322),
            .I(N__25319));
    Span12Mux_v I__3613 (
            .O(N__25319),
            .I(N__25316));
    Odrv12 I__3612 (
            .O(N__25316),
            .I(\current_shift_inst.PI_CTRL.integrator_i_15 ));
    InMux I__3611 (
            .O(N__25313),
            .I(N__25310));
    LocalMux I__3610 (
            .O(N__25310),
            .I(N__25307));
    Odrv12 I__3609 (
            .O(N__25307),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__3608 (
            .O(N__25304),
            .I(bfn_8_18_0_));
    InMux I__3607 (
            .O(N__25301),
            .I(N__25298));
    LocalMux I__3606 (
            .O(N__25298),
            .I(N__25295));
    Odrv4 I__3605 (
            .O(N__25295),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__3604 (
            .O(N__25292),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ));
    InMux I__3603 (
            .O(N__25289),
            .I(N__25286));
    LocalMux I__3602 (
            .O(N__25286),
            .I(N__25283));
    Odrv12 I__3601 (
            .O(N__25283),
            .I(\current_shift_inst.PI_CTRL.integrator_i_17 ));
    CascadeMux I__3600 (
            .O(N__25280),
            .I(N__25277));
    InMux I__3599 (
            .O(N__25277),
            .I(N__25274));
    LocalMux I__3598 (
            .O(N__25274),
            .I(N__25271));
    Odrv4 I__3597 (
            .O(N__25271),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__3596 (
            .O(N__25268),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ));
    InMux I__3595 (
            .O(N__25265),
            .I(N__25262));
    LocalMux I__3594 (
            .O(N__25262),
            .I(N__25259));
    Span4Mux_h I__3593 (
            .O(N__25259),
            .I(N__25256));
    Span4Mux_h I__3592 (
            .O(N__25256),
            .I(N__25253));
    Odrv4 I__3591 (
            .O(N__25253),
            .I(\current_shift_inst.PI_CTRL.integrator_i_18 ));
    InMux I__3590 (
            .O(N__25250),
            .I(N__25247));
    LocalMux I__3589 (
            .O(N__25247),
            .I(N__25244));
    Odrv4 I__3588 (
            .O(N__25244),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__3587 (
            .O(N__25241),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ));
    CascadeMux I__3586 (
            .O(N__25238),
            .I(N__25235));
    InMux I__3585 (
            .O(N__25235),
            .I(N__25232));
    LocalMux I__3584 (
            .O(N__25232),
            .I(N__25229));
    Odrv4 I__3583 (
            .O(N__25229),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__3582 (
            .O(N__25226),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ));
    InMux I__3581 (
            .O(N__25223),
            .I(N__25220));
    LocalMux I__3580 (
            .O(N__25220),
            .I(N__25217));
    Span4Mux_v I__3579 (
            .O(N__25217),
            .I(N__25214));
    Odrv4 I__3578 (
            .O(N__25214),
            .I(\current_shift_inst.PI_CTRL.integrator_i_20 ));
    InMux I__3577 (
            .O(N__25211),
            .I(N__25208));
    LocalMux I__3576 (
            .O(N__25208),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__3575 (
            .O(N__25205),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ));
    InMux I__3574 (
            .O(N__25202),
            .I(N__25199));
    LocalMux I__3573 (
            .O(N__25199),
            .I(\current_shift_inst.PI_CTRL.integrator_i_4 ));
    CascadeMux I__3572 (
            .O(N__25196),
            .I(N__25193));
    InMux I__3571 (
            .O(N__25193),
            .I(N__25190));
    LocalMux I__3570 (
            .O(N__25190),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__3569 (
            .O(N__25187),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ));
    InMux I__3568 (
            .O(N__25184),
            .I(N__25181));
    LocalMux I__3567 (
            .O(N__25181),
            .I(N__25178));
    Odrv4 I__3566 (
            .O(N__25178),
            .I(\current_shift_inst.PI_CTRL.integrator_i_5 ));
    CascadeMux I__3565 (
            .O(N__25175),
            .I(N__25172));
    InMux I__3564 (
            .O(N__25172),
            .I(N__25169));
    LocalMux I__3563 (
            .O(N__25169),
            .I(N__25166));
    Span4Mux_h I__3562 (
            .O(N__25166),
            .I(N__25163));
    Odrv4 I__3561 (
            .O(N__25163),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__3560 (
            .O(N__25160),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ));
    InMux I__3559 (
            .O(N__25157),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ));
    InMux I__3558 (
            .O(N__25154),
            .I(N__25151));
    LocalMux I__3557 (
            .O(N__25151),
            .I(\current_shift_inst.PI_CTRL.integrator_i_7 ));
    CascadeMux I__3556 (
            .O(N__25148),
            .I(N__25145));
    InMux I__3555 (
            .O(N__25145),
            .I(N__25142));
    LocalMux I__3554 (
            .O(N__25142),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11 ));
    CascadeMux I__3553 (
            .O(N__25139),
            .I(N__25136));
    InMux I__3552 (
            .O(N__25136),
            .I(N__25133));
    LocalMux I__3551 (
            .O(N__25133),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__3550 (
            .O(N__25130),
            .I(bfn_8_17_0_));
    InMux I__3549 (
            .O(N__25127),
            .I(N__25124));
    LocalMux I__3548 (
            .O(N__25124),
            .I(N__25121));
    Odrv4 I__3547 (
            .O(N__25121),
            .I(\current_shift_inst.PI_CTRL.integrator_i_8 ));
    InMux I__3546 (
            .O(N__25118),
            .I(N__25115));
    LocalMux I__3545 (
            .O(N__25115),
            .I(N__25112));
    Odrv4 I__3544 (
            .O(N__25112),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__3543 (
            .O(N__25109),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ));
    InMux I__3542 (
            .O(N__25106),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ));
    InMux I__3541 (
            .O(N__25103),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ));
    InMux I__3540 (
            .O(N__25100),
            .I(N__25097));
    LocalMux I__3539 (
            .O(N__25097),
            .I(N__25094));
    Odrv4 I__3538 (
            .O(N__25094),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__3537 (
            .O(N__25091),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ));
    InMux I__3536 (
            .O(N__25088),
            .I(N__25085));
    LocalMux I__3535 (
            .O(N__25085),
            .I(N__25082));
    Odrv12 I__3534 (
            .O(N__25082),
            .I(\current_shift_inst.PI_CTRL.integrator_i_12 ));
    InMux I__3533 (
            .O(N__25079),
            .I(N__25076));
    LocalMux I__3532 (
            .O(N__25076),
            .I(N__25073));
    Span4Mux_v I__3531 (
            .O(N__25073),
            .I(N__25070));
    Odrv4 I__3530 (
            .O(N__25070),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__3529 (
            .O(N__25067),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ));
    InMux I__3528 (
            .O(N__25064),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ));
    InMux I__3527 (
            .O(N__25061),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ));
    InMux I__3526 (
            .O(N__25058),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ));
    InMux I__3525 (
            .O(N__25055),
            .I(N__25052));
    LocalMux I__3524 (
            .O(N__25052),
            .I(N__25049));
    Odrv4 I__3523 (
            .O(N__25049),
            .I(\current_shift_inst.PI_CTRL.integrator_i_3 ));
    CascadeMux I__3522 (
            .O(N__25046),
            .I(N__25043));
    InMux I__3521 (
            .O(N__25043),
            .I(N__25040));
    LocalMux I__3520 (
            .O(N__25040),
            .I(N__25037));
    Span4Mux_v I__3519 (
            .O(N__25037),
            .I(N__25034));
    Odrv4 I__3518 (
            .O(N__25034),
            .I(\current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7 ));
    InMux I__3517 (
            .O(N__25031),
            .I(N__25028));
    LocalMux I__3516 (
            .O(N__25028),
            .I(N__25025));
    Odrv4 I__3515 (
            .O(N__25025),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__3514 (
            .O(N__25022),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ));
    CascadeMux I__3513 (
            .O(N__25019),
            .I(N__25015));
    InMux I__3512 (
            .O(N__25018),
            .I(N__25012));
    InMux I__3511 (
            .O(N__25015),
            .I(N__25009));
    LocalMux I__3510 (
            .O(N__25012),
            .I(N__25005));
    LocalMux I__3509 (
            .O(N__25009),
            .I(N__25002));
    InMux I__3508 (
            .O(N__25008),
            .I(N__24999));
    Span4Mux_h I__3507 (
            .O(N__25005),
            .I(N__24994));
    Span4Mux_h I__3506 (
            .O(N__25002),
            .I(N__24994));
    LocalMux I__3505 (
            .O(N__24999),
            .I(N__24989));
    Span4Mux_h I__3504 (
            .O(N__24994),
            .I(N__24986));
    InMux I__3503 (
            .O(N__24993),
            .I(N__24981));
    InMux I__3502 (
            .O(N__24992),
            .I(N__24981));
    Odrv4 I__3501 (
            .O(N__24989),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__3500 (
            .O(N__24986),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__3499 (
            .O(N__24981),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__3498 (
            .O(N__24974),
            .I(N__24971));
    LocalMux I__3497 (
            .O(N__24971),
            .I(N__24968));
    Odrv4 I__3496 (
            .O(N__24968),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt24 ));
    InMux I__3495 (
            .O(N__24965),
            .I(N__24959));
    InMux I__3494 (
            .O(N__24964),
            .I(N__24959));
    LocalMux I__3493 (
            .O(N__24959),
            .I(N__24956));
    Odrv4 I__3492 (
            .O(N__24956),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    InMux I__3491 (
            .O(N__24953),
            .I(N__24948));
    InMux I__3490 (
            .O(N__24952),
            .I(N__24943));
    InMux I__3489 (
            .O(N__24951),
            .I(N__24943));
    LocalMux I__3488 (
            .O(N__24948),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    LocalMux I__3487 (
            .O(N__24943),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    CascadeMux I__3486 (
            .O(N__24938),
            .I(N__24935));
    InMux I__3485 (
            .O(N__24935),
            .I(N__24928));
    InMux I__3484 (
            .O(N__24934),
            .I(N__24928));
    InMux I__3483 (
            .O(N__24933),
            .I(N__24925));
    LocalMux I__3482 (
            .O(N__24928),
            .I(N__24922));
    LocalMux I__3481 (
            .O(N__24925),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__3480 (
            .O(N__24922),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    CascadeMux I__3479 (
            .O(N__24917),
            .I(N__24914));
    InMux I__3478 (
            .O(N__24914),
            .I(N__24911));
    LocalMux I__3477 (
            .O(N__24911),
            .I(N__24908));
    Odrv4 I__3476 (
            .O(N__24908),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ));
    CascadeMux I__3475 (
            .O(N__24905),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_));
    InMux I__3474 (
            .O(N__24902),
            .I(N__24899));
    LocalMux I__3473 (
            .O(N__24899),
            .I(N__24896));
    Odrv4 I__3472 (
            .O(N__24896),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ));
    InMux I__3471 (
            .O(N__24893),
            .I(N__24886));
    InMux I__3470 (
            .O(N__24892),
            .I(N__24886));
    InMux I__3469 (
            .O(N__24891),
            .I(N__24883));
    LocalMux I__3468 (
            .O(N__24886),
            .I(N__24880));
    LocalMux I__3467 (
            .O(N__24883),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv4 I__3466 (
            .O(N__24880),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    CascadeMux I__3465 (
            .O(N__24875),
            .I(N__24872));
    InMux I__3464 (
            .O(N__24872),
            .I(N__24865));
    InMux I__3463 (
            .O(N__24871),
            .I(N__24865));
    InMux I__3462 (
            .O(N__24870),
            .I(N__24862));
    LocalMux I__3461 (
            .O(N__24865),
            .I(N__24859));
    LocalMux I__3460 (
            .O(N__24862),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__3459 (
            .O(N__24859),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__3458 (
            .O(N__24854),
            .I(N__24848));
    InMux I__3457 (
            .O(N__24853),
            .I(N__24848));
    LocalMux I__3456 (
            .O(N__24848),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ));
    CascadeMux I__3455 (
            .O(N__24845),
            .I(N__24842));
    InMux I__3454 (
            .O(N__24842),
            .I(N__24839));
    LocalMux I__3453 (
            .O(N__24839),
            .I(N__24836));
    Span4Mux_h I__3452 (
            .O(N__24836),
            .I(N__24833));
    Odrv4 I__3451 (
            .O(N__24833),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt26 ));
    CascadeMux I__3450 (
            .O(N__24830),
            .I(N__24827));
    InMux I__3449 (
            .O(N__24827),
            .I(N__24821));
    InMux I__3448 (
            .O(N__24826),
            .I(N__24821));
    LocalMux I__3447 (
            .O(N__24821),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    CascadeMux I__3446 (
            .O(N__24818),
            .I(N__24815));
    InMux I__3445 (
            .O(N__24815),
            .I(N__24809));
    InMux I__3444 (
            .O(N__24814),
            .I(N__24809));
    LocalMux I__3443 (
            .O(N__24809),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    CEMux I__3442 (
            .O(N__24806),
            .I(N__24785));
    CEMux I__3441 (
            .O(N__24805),
            .I(N__24785));
    CEMux I__3440 (
            .O(N__24804),
            .I(N__24785));
    CEMux I__3439 (
            .O(N__24803),
            .I(N__24785));
    CEMux I__3438 (
            .O(N__24802),
            .I(N__24785));
    CEMux I__3437 (
            .O(N__24801),
            .I(N__24785));
    CEMux I__3436 (
            .O(N__24800),
            .I(N__24785));
    GlobalMux I__3435 (
            .O(N__24785),
            .I(N__24782));
    gio2CtrlBuf I__3434 (
            .O(N__24782),
            .I(\phase_controller_inst2.stoper_tr.un1_start_g ));
    CascadeMux I__3433 (
            .O(N__24779),
            .I(\phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_ ));
    InMux I__3432 (
            .O(N__24776),
            .I(N__24770));
    InMux I__3431 (
            .O(N__24775),
            .I(N__24770));
    LocalMux I__3430 (
            .O(N__24770),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__3429 (
            .O(N__24767),
            .I(N__24764));
    LocalMux I__3428 (
            .O(N__24764),
            .I(N__24761));
    Odrv4 I__3427 (
            .O(N__24761),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df30 ));
    CascadeMux I__3426 (
            .O(N__24758),
            .I(N__24755));
    InMux I__3425 (
            .O(N__24755),
            .I(N__24751));
    InMux I__3424 (
            .O(N__24754),
            .I(N__24748));
    LocalMux I__3423 (
            .O(N__24751),
            .I(N__24745));
    LocalMux I__3422 (
            .O(N__24748),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    Odrv4 I__3421 (
            .O(N__24745),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    InMux I__3420 (
            .O(N__24740),
            .I(N__24737));
    LocalMux I__3419 (
            .O(N__24737),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ));
    CascadeMux I__3418 (
            .O(N__24734),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__3417 (
            .O(N__24731),
            .I(N__24728));
    InMux I__3416 (
            .O(N__24728),
            .I(N__24725));
    LocalMux I__3415 (
            .O(N__24725),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    InMux I__3414 (
            .O(N__24722),
            .I(N__24719));
    LocalMux I__3413 (
            .O(N__24719),
            .I(N__24715));
    InMux I__3412 (
            .O(N__24718),
            .I(N__24710));
    Span4Mux_h I__3411 (
            .O(N__24715),
            .I(N__24707));
    InMux I__3410 (
            .O(N__24714),
            .I(N__24702));
    InMux I__3409 (
            .O(N__24713),
            .I(N__24702));
    LocalMux I__3408 (
            .O(N__24710),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__3407 (
            .O(N__24707),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__3406 (
            .O(N__24702),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__3405 (
            .O(N__24695),
            .I(N__24692));
    LocalMux I__3404 (
            .O(N__24692),
            .I(N__24689));
    Span4Mux_v I__3403 (
            .O(N__24689),
            .I(N__24685));
    InMux I__3402 (
            .O(N__24688),
            .I(N__24682));
    Odrv4 I__3401 (
            .O(N__24685),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__3400 (
            .O(N__24682),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__3399 (
            .O(N__24677),
            .I(N__24674));
    InMux I__3398 (
            .O(N__24674),
            .I(N__24671));
    LocalMux I__3397 (
            .O(N__24671),
            .I(N__24668));
    Odrv4 I__3396 (
            .O(N__24668),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ));
    CascadeMux I__3395 (
            .O(N__24665),
            .I(N__24661));
    CascadeMux I__3394 (
            .O(N__24664),
            .I(N__24657));
    InMux I__3393 (
            .O(N__24661),
            .I(N__24650));
    InMux I__3392 (
            .O(N__24660),
            .I(N__24650));
    InMux I__3391 (
            .O(N__24657),
            .I(N__24650));
    LocalMux I__3390 (
            .O(N__24650),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    InMux I__3389 (
            .O(N__24647),
            .I(N__24644));
    LocalMux I__3388 (
            .O(N__24644),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__3387 (
            .O(N__24641),
            .I(N__24638));
    InMux I__3386 (
            .O(N__24638),
            .I(N__24635));
    LocalMux I__3385 (
            .O(N__24635),
            .I(N__24632));
    Odrv4 I__3384 (
            .O(N__24632),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt22 ));
    InMux I__3383 (
            .O(N__24629),
            .I(N__24622));
    InMux I__3382 (
            .O(N__24628),
            .I(N__24622));
    InMux I__3381 (
            .O(N__24627),
            .I(N__24619));
    LocalMux I__3380 (
            .O(N__24622),
            .I(N__24616));
    LocalMux I__3379 (
            .O(N__24619),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__3378 (
            .O(N__24616),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    CascadeMux I__3377 (
            .O(N__24611),
            .I(N__24608));
    InMux I__3376 (
            .O(N__24608),
            .I(N__24602));
    InMux I__3375 (
            .O(N__24607),
            .I(N__24602));
    LocalMux I__3374 (
            .O(N__24602),
            .I(N__24598));
    InMux I__3373 (
            .O(N__24601),
            .I(N__24595));
    Span4Mux_h I__3372 (
            .O(N__24598),
            .I(N__24592));
    LocalMux I__3371 (
            .O(N__24595),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__3370 (
            .O(N__24592),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__3369 (
            .O(N__24587),
            .I(N__24584));
    LocalMux I__3368 (
            .O(N__24584),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ));
    InMux I__3367 (
            .O(N__24581),
            .I(N__24575));
    InMux I__3366 (
            .O(N__24580),
            .I(N__24575));
    LocalMux I__3365 (
            .O(N__24575),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ));
    CascadeMux I__3364 (
            .O(N__24572),
            .I(N__24569));
    InMux I__3363 (
            .O(N__24569),
            .I(N__24563));
    InMux I__3362 (
            .O(N__24568),
            .I(N__24563));
    LocalMux I__3361 (
            .O(N__24563),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ));
    CascadeMux I__3360 (
            .O(N__24560),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12_cascade_));
    InMux I__3359 (
            .O(N__24557),
            .I(N__24554));
    LocalMux I__3358 (
            .O(N__24554),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__3357 (
            .O(N__24551),
            .I(N__24548));
    InMux I__3356 (
            .O(N__24548),
            .I(N__24545));
    LocalMux I__3355 (
            .O(N__24545),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__3354 (
            .O(N__24542),
            .I(N__24539));
    InMux I__3353 (
            .O(N__24539),
            .I(N__24536));
    LocalMux I__3352 (
            .O(N__24536),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    InMux I__3351 (
            .O(N__24533),
            .I(N__24530));
    LocalMux I__3350 (
            .O(N__24530),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    InMux I__3349 (
            .O(N__24527),
            .I(N__24524));
    LocalMux I__3348 (
            .O(N__24524),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    InMux I__3347 (
            .O(N__24521),
            .I(N__24518));
    LocalMux I__3346 (
            .O(N__24518),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    InMux I__3345 (
            .O(N__24515),
            .I(N__24506));
    InMux I__3344 (
            .O(N__24514),
            .I(N__24506));
    InMux I__3343 (
            .O(N__24513),
            .I(N__24506));
    LocalMux I__3342 (
            .O(N__24506),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    CascadeMux I__3341 (
            .O(N__24503),
            .I(N__24498));
    InMux I__3340 (
            .O(N__24502),
            .I(N__24491));
    InMux I__3339 (
            .O(N__24501),
            .I(N__24491));
    InMux I__3338 (
            .O(N__24498),
            .I(N__24491));
    LocalMux I__3337 (
            .O(N__24491),
            .I(N__24487));
    InMux I__3336 (
            .O(N__24490),
            .I(N__24484));
    Span4Mux_v I__3335 (
            .O(N__24487),
            .I(N__24481));
    LocalMux I__3334 (
            .O(N__24484),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__3333 (
            .O(N__24481),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__3332 (
            .O(N__24476),
            .I(N__24467));
    InMux I__3331 (
            .O(N__24475),
            .I(N__24467));
    InMux I__3330 (
            .O(N__24474),
            .I(N__24467));
    LocalMux I__3329 (
            .O(N__24467),
            .I(N__24463));
    InMux I__3328 (
            .O(N__24466),
            .I(N__24460));
    Span4Mux_v I__3327 (
            .O(N__24463),
            .I(N__24457));
    LocalMux I__3326 (
            .O(N__24460),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__3325 (
            .O(N__24457),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    CascadeMux I__3324 (
            .O(N__24452),
            .I(N__24449));
    InMux I__3323 (
            .O(N__24449),
            .I(N__24446));
    LocalMux I__3322 (
            .O(N__24446),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    CascadeMux I__3321 (
            .O(N__24443),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_));
    InMux I__3320 (
            .O(N__24440),
            .I(N__24437));
    LocalMux I__3319 (
            .O(N__24437),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    InMux I__3318 (
            .O(N__24434),
            .I(N__24428));
    InMux I__3317 (
            .O(N__24433),
            .I(N__24428));
    LocalMux I__3316 (
            .O(N__24428),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    InMux I__3315 (
            .O(N__24425),
            .I(N__24422));
    LocalMux I__3314 (
            .O(N__24422),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__3313 (
            .O(N__24419),
            .I(N__24416));
    InMux I__3312 (
            .O(N__24416),
            .I(N__24410));
    InMux I__3311 (
            .O(N__24415),
            .I(N__24410));
    LocalMux I__3310 (
            .O(N__24410),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    InMux I__3309 (
            .O(N__24407),
            .I(N__24404));
    LocalMux I__3308 (
            .O(N__24404),
            .I(N__24401));
    Odrv4 I__3307 (
            .O(N__24401),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__3306 (
            .O(N__24398),
            .I(N__24395));
    InMux I__3305 (
            .O(N__24395),
            .I(N__24392));
    LocalMux I__3304 (
            .O(N__24392),
            .I(N__24389));
    Odrv4 I__3303 (
            .O(N__24389),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__3302 (
            .O(N__24386),
            .I(N__24383));
    InMux I__3301 (
            .O(N__24383),
            .I(N__24380));
    LocalMux I__3300 (
            .O(N__24380),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    InMux I__3299 (
            .O(N__24377),
            .I(N__24371));
    InMux I__3298 (
            .O(N__24376),
            .I(N__24371));
    LocalMux I__3297 (
            .O(N__24371),
            .I(N__24367));
    InMux I__3296 (
            .O(N__24370),
            .I(N__24364));
    Span4Mux_v I__3295 (
            .O(N__24367),
            .I(N__24361));
    LocalMux I__3294 (
            .O(N__24364),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__3293 (
            .O(N__24361),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__3292 (
            .O(N__24356),
            .I(N__24353));
    InMux I__3291 (
            .O(N__24353),
            .I(N__24347));
    InMux I__3290 (
            .O(N__24352),
            .I(N__24347));
    LocalMux I__3289 (
            .O(N__24347),
            .I(N__24344));
    Span4Mux_v I__3288 (
            .O(N__24344),
            .I(N__24340));
    InMux I__3287 (
            .O(N__24343),
            .I(N__24337));
    Span4Mux_h I__3286 (
            .O(N__24340),
            .I(N__24334));
    LocalMux I__3285 (
            .O(N__24337),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__3284 (
            .O(N__24334),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__3283 (
            .O(N__24329),
            .I(N__24326));
    LocalMux I__3282 (
            .O(N__24326),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    InMux I__3281 (
            .O(N__24323),
            .I(N__24317));
    InMux I__3280 (
            .O(N__24322),
            .I(N__24317));
    LocalMux I__3279 (
            .O(N__24317),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__3278 (
            .O(N__24314),
            .I(N__24311));
    InMux I__3277 (
            .O(N__24311),
            .I(N__24305));
    InMux I__3276 (
            .O(N__24310),
            .I(N__24305));
    LocalMux I__3275 (
            .O(N__24305),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__3274 (
            .O(N__24302),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ));
    CascadeMux I__3273 (
            .O(N__24299),
            .I(N__24296));
    InMux I__3272 (
            .O(N__24296),
            .I(N__24293));
    LocalMux I__3271 (
            .O(N__24293),
            .I(N__24290));
    Span4Mux_v I__3270 (
            .O(N__24290),
            .I(N__24287));
    Odrv4 I__3269 (
            .O(N__24287),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt20 ));
    InMux I__3268 (
            .O(N__24284),
            .I(N__24278));
    InMux I__3267 (
            .O(N__24283),
            .I(N__24278));
    LocalMux I__3266 (
            .O(N__24278),
            .I(N__24274));
    InMux I__3265 (
            .O(N__24277),
            .I(N__24271));
    Span4Mux_v I__3264 (
            .O(N__24274),
            .I(N__24268));
    LocalMux I__3263 (
            .O(N__24271),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__3262 (
            .O(N__24268),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    CascadeMux I__3261 (
            .O(N__24263),
            .I(N__24260));
    InMux I__3260 (
            .O(N__24260),
            .I(N__24254));
    InMux I__3259 (
            .O(N__24259),
            .I(N__24254));
    LocalMux I__3258 (
            .O(N__24254),
            .I(N__24250));
    InMux I__3257 (
            .O(N__24253),
            .I(N__24247));
    Span4Mux_v I__3256 (
            .O(N__24250),
            .I(N__24244));
    LocalMux I__3255 (
            .O(N__24247),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__3254 (
            .O(N__24244),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__3253 (
            .O(N__24239),
            .I(N__24236));
    LocalMux I__3252 (
            .O(N__24236),
            .I(N__24233));
    Span4Mux_v I__3251 (
            .O(N__24233),
            .I(N__24230));
    Odrv4 I__3250 (
            .O(N__24230),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ));
    InMux I__3249 (
            .O(N__24227),
            .I(N__24221));
    InMux I__3248 (
            .O(N__24226),
            .I(N__24214));
    InMux I__3247 (
            .O(N__24225),
            .I(N__24214));
    InMux I__3246 (
            .O(N__24224),
            .I(N__24214));
    LocalMux I__3245 (
            .O(N__24221),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__3244 (
            .O(N__24214),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    CascadeMux I__3243 (
            .O(N__24209),
            .I(N__24206));
    InMux I__3242 (
            .O(N__24206),
            .I(N__24201));
    InMux I__3241 (
            .O(N__24205),
            .I(N__24198));
    InMux I__3240 (
            .O(N__24204),
            .I(N__24195));
    LocalMux I__3239 (
            .O(N__24201),
            .I(N__24190));
    LocalMux I__3238 (
            .O(N__24198),
            .I(N__24190));
    LocalMux I__3237 (
            .O(N__24195),
            .I(N__24183));
    Span4Mux_h I__3236 (
            .O(N__24190),
            .I(N__24183));
    InMux I__3235 (
            .O(N__24189),
            .I(N__24178));
    InMux I__3234 (
            .O(N__24188),
            .I(N__24178));
    Odrv4 I__3233 (
            .O(N__24183),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__3232 (
            .O(N__24178),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__3231 (
            .O(N__24173),
            .I(N__24170));
    LocalMux I__3230 (
            .O(N__24170),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__3229 (
            .O(N__24167),
            .I(N__24164));
    LocalMux I__3228 (
            .O(N__24164),
            .I(N__24161));
    Odrv12 I__3227 (
            .O(N__24161),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ));
    CascadeMux I__3226 (
            .O(N__24158),
            .I(N__24155));
    InMux I__3225 (
            .O(N__24155),
            .I(N__24152));
    LocalMux I__3224 (
            .O(N__24152),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    InMux I__3223 (
            .O(N__24149),
            .I(N__24146));
    LocalMux I__3222 (
            .O(N__24146),
            .I(N__24143));
    Odrv12 I__3221 (
            .O(N__24143),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ));
    InMux I__3220 (
            .O(N__24140),
            .I(N__24137));
    LocalMux I__3219 (
            .O(N__24137),
            .I(N__24134));
    Odrv12 I__3218 (
            .O(N__24134),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    CascadeMux I__3217 (
            .O(N__24131),
            .I(N__24127));
    InMux I__3216 (
            .O(N__24130),
            .I(N__24122));
    InMux I__3215 (
            .O(N__24127),
            .I(N__24122));
    LocalMux I__3214 (
            .O(N__24122),
            .I(N__24118));
    InMux I__3213 (
            .O(N__24121),
            .I(N__24115));
    Span4Mux_h I__3212 (
            .O(N__24118),
            .I(N__24112));
    LocalMux I__3211 (
            .O(N__24115),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__3210 (
            .O(N__24112),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__3209 (
            .O(N__24107),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__3208 (
            .O(N__24104),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__3207 (
            .O(N__24101),
            .I(N__24078));
    InMux I__3206 (
            .O(N__24100),
            .I(N__24078));
    InMux I__3205 (
            .O(N__24099),
            .I(N__24078));
    InMux I__3204 (
            .O(N__24098),
            .I(N__24078));
    InMux I__3203 (
            .O(N__24097),
            .I(N__24071));
    InMux I__3202 (
            .O(N__24096),
            .I(N__24071));
    InMux I__3201 (
            .O(N__24095),
            .I(N__24071));
    InMux I__3200 (
            .O(N__24094),
            .I(N__24062));
    InMux I__3199 (
            .O(N__24093),
            .I(N__24062));
    InMux I__3198 (
            .O(N__24092),
            .I(N__24062));
    InMux I__3197 (
            .O(N__24091),
            .I(N__24062));
    InMux I__3196 (
            .O(N__24090),
            .I(N__24053));
    InMux I__3195 (
            .O(N__24089),
            .I(N__24053));
    InMux I__3194 (
            .O(N__24088),
            .I(N__24053));
    InMux I__3193 (
            .O(N__24087),
            .I(N__24053));
    LocalMux I__3192 (
            .O(N__24078),
            .I(N__24034));
    LocalMux I__3191 (
            .O(N__24071),
            .I(N__24027));
    LocalMux I__3190 (
            .O(N__24062),
            .I(N__24027));
    LocalMux I__3189 (
            .O(N__24053),
            .I(N__24027));
    InMux I__3188 (
            .O(N__24052),
            .I(N__24020));
    InMux I__3187 (
            .O(N__24051),
            .I(N__24020));
    InMux I__3186 (
            .O(N__24050),
            .I(N__24020));
    InMux I__3185 (
            .O(N__24049),
            .I(N__24011));
    InMux I__3184 (
            .O(N__24048),
            .I(N__24011));
    InMux I__3183 (
            .O(N__24047),
            .I(N__24011));
    InMux I__3182 (
            .O(N__24046),
            .I(N__24011));
    InMux I__3181 (
            .O(N__24045),
            .I(N__24002));
    InMux I__3180 (
            .O(N__24044),
            .I(N__24002));
    InMux I__3179 (
            .O(N__24043),
            .I(N__24002));
    InMux I__3178 (
            .O(N__24042),
            .I(N__24002));
    InMux I__3177 (
            .O(N__24041),
            .I(N__23993));
    InMux I__3176 (
            .O(N__24040),
            .I(N__23993));
    InMux I__3175 (
            .O(N__24039),
            .I(N__23993));
    InMux I__3174 (
            .O(N__24038),
            .I(N__23993));
    IoInMux I__3173 (
            .O(N__24037),
            .I(N__23990));
    Span4Mux_v I__3172 (
            .O(N__24034),
            .I(N__23977));
    Span4Mux_v I__3171 (
            .O(N__24027),
            .I(N__23977));
    LocalMux I__3170 (
            .O(N__24020),
            .I(N__23977));
    LocalMux I__3169 (
            .O(N__24011),
            .I(N__23977));
    LocalMux I__3168 (
            .O(N__24002),
            .I(N__23977));
    LocalMux I__3167 (
            .O(N__23993),
            .I(N__23977));
    LocalMux I__3166 (
            .O(N__23990),
            .I(N__23974));
    Span4Mux_v I__3165 (
            .O(N__23977),
            .I(N__23971));
    Span12Mux_s8_v I__3164 (
            .O(N__23974),
            .I(N__23968));
    Odrv4 I__3163 (
            .O(N__23971),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv12 I__3162 (
            .O(N__23968),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__3161 (
            .O(N__23963),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__3160 (
            .O(N__23960),
            .I(N__23957));
    LocalMux I__3159 (
            .O(N__23957),
            .I(N__23954));
    Odrv4 I__3158 (
            .O(N__23954),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__3157 (
            .O(N__23951),
            .I(N__23948));
    LocalMux I__3156 (
            .O(N__23948),
            .I(N__23945));
    Span4Mux_v I__3155 (
            .O(N__23945),
            .I(N__23942));
    Odrv4 I__3154 (
            .O(N__23942),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    CascadeMux I__3153 (
            .O(N__23939),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    CascadeMux I__3152 (
            .O(N__23936),
            .I(\current_shift_inst.PI_CTRL.N_72_cascade_ ));
    InMux I__3151 (
            .O(N__23933),
            .I(N__23930));
    LocalMux I__3150 (
            .O(N__23930),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    InMux I__3149 (
            .O(N__23927),
            .I(N__23924));
    LocalMux I__3148 (
            .O(N__23924),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    InMux I__3147 (
            .O(N__23921),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__3146 (
            .O(N__23918),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__3145 (
            .O(N__23915),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__3144 (
            .O(N__23912),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__3143 (
            .O(N__23909),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__3142 (
            .O(N__23906),
            .I(bfn_7_15_0_));
    InMux I__3141 (
            .O(N__23903),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__3140 (
            .O(N__23900),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    CascadeMux I__3139 (
            .O(N__23897),
            .I(N__23894));
    InMux I__3138 (
            .O(N__23894),
            .I(N__23890));
    InMux I__3137 (
            .O(N__23893),
            .I(N__23887));
    LocalMux I__3136 (
            .O(N__23890),
            .I(N__23881));
    LocalMux I__3135 (
            .O(N__23887),
            .I(N__23881));
    InMux I__3134 (
            .O(N__23886),
            .I(N__23878));
    Span4Mux_h I__3133 (
            .O(N__23881),
            .I(N__23875));
    LocalMux I__3132 (
            .O(N__23878),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__3131 (
            .O(N__23875),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__3130 (
            .O(N__23870),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__3129 (
            .O(N__23867),
            .I(N__23863));
    InMux I__3128 (
            .O(N__23866),
            .I(N__23860));
    LocalMux I__3127 (
            .O(N__23863),
            .I(N__23857));
    LocalMux I__3126 (
            .O(N__23860),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__3125 (
            .O(N__23857),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__3124 (
            .O(N__23852),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__3123 (
            .O(N__23849),
            .I(N__23845));
    InMux I__3122 (
            .O(N__23848),
            .I(N__23842));
    LocalMux I__3121 (
            .O(N__23845),
            .I(N__23839));
    LocalMux I__3120 (
            .O(N__23842),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__3119 (
            .O(N__23839),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__3118 (
            .O(N__23834),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__3117 (
            .O(N__23831),
            .I(N__23828));
    LocalMux I__3116 (
            .O(N__23828),
            .I(N__23824));
    InMux I__3115 (
            .O(N__23827),
            .I(N__23821));
    Span4Mux_v I__3114 (
            .O(N__23824),
            .I(N__23818));
    LocalMux I__3113 (
            .O(N__23821),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__3112 (
            .O(N__23818),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__3111 (
            .O(N__23813),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__3110 (
            .O(N__23810),
            .I(N__23806));
    InMux I__3109 (
            .O(N__23809),
            .I(N__23803));
    LocalMux I__3108 (
            .O(N__23806),
            .I(N__23800));
    LocalMux I__3107 (
            .O(N__23803),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__3106 (
            .O(N__23800),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__3105 (
            .O(N__23795),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__3104 (
            .O(N__23792),
            .I(N__23788));
    InMux I__3103 (
            .O(N__23791),
            .I(N__23785));
    LocalMux I__3102 (
            .O(N__23788),
            .I(N__23782));
    LocalMux I__3101 (
            .O(N__23785),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv12 I__3100 (
            .O(N__23782),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__3099 (
            .O(N__23777),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__3098 (
            .O(N__23774),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__3097 (
            .O(N__23771),
            .I(bfn_7_14_0_));
    InMux I__3096 (
            .O(N__23768),
            .I(N__23761));
    InMux I__3095 (
            .O(N__23767),
            .I(N__23761));
    InMux I__3094 (
            .O(N__23766),
            .I(N__23758));
    LocalMux I__3093 (
            .O(N__23761),
            .I(N__23755));
    LocalMux I__3092 (
            .O(N__23758),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv12 I__3091 (
            .O(N__23755),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__3090 (
            .O(N__23750),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    CascadeMux I__3089 (
            .O(N__23747),
            .I(N__23744));
    InMux I__3088 (
            .O(N__23744),
            .I(N__23738));
    InMux I__3087 (
            .O(N__23743),
            .I(N__23738));
    LocalMux I__3086 (
            .O(N__23738),
            .I(N__23734));
    InMux I__3085 (
            .O(N__23737),
            .I(N__23731));
    Span4Mux_v I__3084 (
            .O(N__23734),
            .I(N__23728));
    LocalMux I__3083 (
            .O(N__23731),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__3082 (
            .O(N__23728),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__3081 (
            .O(N__23723),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__3080 (
            .O(N__23720),
            .I(N__23716));
    InMux I__3079 (
            .O(N__23719),
            .I(N__23713));
    LocalMux I__3078 (
            .O(N__23716),
            .I(N__23710));
    LocalMux I__3077 (
            .O(N__23713),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__3076 (
            .O(N__23710),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__3075 (
            .O(N__23705),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__3074 (
            .O(N__23702),
            .I(N__23698));
    InMux I__3073 (
            .O(N__23701),
            .I(N__23695));
    LocalMux I__3072 (
            .O(N__23698),
            .I(N__23692));
    LocalMux I__3071 (
            .O(N__23695),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__3070 (
            .O(N__23692),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__3069 (
            .O(N__23687),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__3068 (
            .O(N__23684),
            .I(N__23681));
    LocalMux I__3067 (
            .O(N__23681),
            .I(N__23677));
    InMux I__3066 (
            .O(N__23680),
            .I(N__23674));
    Span4Mux_v I__3065 (
            .O(N__23677),
            .I(N__23671));
    LocalMux I__3064 (
            .O(N__23674),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__3063 (
            .O(N__23671),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__3062 (
            .O(N__23666),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__3061 (
            .O(N__23663),
            .I(N__23660));
    LocalMux I__3060 (
            .O(N__23660),
            .I(N__23656));
    InMux I__3059 (
            .O(N__23659),
            .I(N__23653));
    Span4Mux_v I__3058 (
            .O(N__23656),
            .I(N__23650));
    LocalMux I__3057 (
            .O(N__23653),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__3056 (
            .O(N__23650),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__3055 (
            .O(N__23645),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__3054 (
            .O(N__23642),
            .I(N__23638));
    InMux I__3053 (
            .O(N__23641),
            .I(N__23635));
    LocalMux I__3052 (
            .O(N__23638),
            .I(N__23632));
    LocalMux I__3051 (
            .O(N__23635),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__3050 (
            .O(N__23632),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__3049 (
            .O(N__23627),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__3048 (
            .O(N__23624),
            .I(N__23620));
    InMux I__3047 (
            .O(N__23623),
            .I(N__23617));
    LocalMux I__3046 (
            .O(N__23620),
            .I(N__23614));
    LocalMux I__3045 (
            .O(N__23617),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv12 I__3044 (
            .O(N__23614),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__3043 (
            .O(N__23609),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__3042 (
            .O(N__23606),
            .I(N__23603));
    LocalMux I__3041 (
            .O(N__23603),
            .I(N__23599));
    InMux I__3040 (
            .O(N__23602),
            .I(N__23596));
    Span4Mux_h I__3039 (
            .O(N__23599),
            .I(N__23593));
    LocalMux I__3038 (
            .O(N__23596),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__3037 (
            .O(N__23593),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__3036 (
            .O(N__23588),
            .I(bfn_7_13_0_));
    InMux I__3035 (
            .O(N__23585),
            .I(N__23582));
    LocalMux I__3034 (
            .O(N__23582),
            .I(N__23578));
    InMux I__3033 (
            .O(N__23581),
            .I(N__23575));
    Span4Mux_h I__3032 (
            .O(N__23578),
            .I(N__23572));
    LocalMux I__3031 (
            .O(N__23575),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__3030 (
            .O(N__23572),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__3029 (
            .O(N__23567),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__3028 (
            .O(N__23564),
            .I(N__23561));
    LocalMux I__3027 (
            .O(N__23561),
            .I(N__23558));
    Odrv4 I__3026 (
            .O(N__23558),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ));
    CascadeMux I__3025 (
            .O(N__23555),
            .I(N__23552));
    InMux I__3024 (
            .O(N__23552),
            .I(N__23549));
    LocalMux I__3023 (
            .O(N__23549),
            .I(N__23546));
    Odrv4 I__3022 (
            .O(N__23546),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt28 ));
    InMux I__3021 (
            .O(N__23543),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ));
    InMux I__3020 (
            .O(N__23540),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    InMux I__3019 (
            .O(N__23537),
            .I(N__23534));
    LocalMux I__3018 (
            .O(N__23534),
            .I(N__23529));
    InMux I__3017 (
            .O(N__23533),
            .I(N__23526));
    InMux I__3016 (
            .O(N__23532),
            .I(N__23523));
    Span4Mux_v I__3015 (
            .O(N__23529),
            .I(N__23518));
    LocalMux I__3014 (
            .O(N__23526),
            .I(N__23518));
    LocalMux I__3013 (
            .O(N__23523),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__3012 (
            .O(N__23518),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__3011 (
            .O(N__23513),
            .I(N__23509));
    InMux I__3010 (
            .O(N__23512),
            .I(N__23506));
    LocalMux I__3009 (
            .O(N__23509),
            .I(N__23503));
    LocalMux I__3008 (
            .O(N__23506),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__3007 (
            .O(N__23503),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__3006 (
            .O(N__23498),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__3005 (
            .O(N__23495),
            .I(N__23492));
    InMux I__3004 (
            .O(N__23492),
            .I(N__23489));
    LocalMux I__3003 (
            .O(N__23489),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__3002 (
            .O(N__23486),
            .I(N__23483));
    LocalMux I__3001 (
            .O(N__23483),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__3000 (
            .O(N__23480),
            .I(N__23477));
    LocalMux I__2999 (
            .O(N__23477),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__2998 (
            .O(N__23474),
            .I(N__23471));
    InMux I__2997 (
            .O(N__23471),
            .I(N__23468));
    LocalMux I__2996 (
            .O(N__23468),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__2995 (
            .O(N__23465),
            .I(N__23462));
    InMux I__2994 (
            .O(N__23462),
            .I(N__23459));
    LocalMux I__2993 (
            .O(N__23459),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__2992 (
            .O(N__23456),
            .I(N__23453));
    InMux I__2991 (
            .O(N__23453),
            .I(N__23450));
    LocalMux I__2990 (
            .O(N__23450),
            .I(N__23447));
    Odrv4 I__2989 (
            .O(N__23447),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__2988 (
            .O(N__23444),
            .I(N__23441));
    LocalMux I__2987 (
            .O(N__23441),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__2986 (
            .O(N__23438),
            .I(N__23435));
    LocalMux I__2985 (
            .O(N__23435),
            .I(N__23432));
    Odrv12 I__2984 (
            .O(N__23432),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    CascadeMux I__2983 (
            .O(N__23429),
            .I(N__23426));
    InMux I__2982 (
            .O(N__23426),
            .I(N__23423));
    LocalMux I__2981 (
            .O(N__23423),
            .I(N__23420));
    Odrv12 I__2980 (
            .O(N__23420),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    CascadeMux I__2979 (
            .O(N__23417),
            .I(N__23414));
    InMux I__2978 (
            .O(N__23414),
            .I(N__23411));
    LocalMux I__2977 (
            .O(N__23411),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__2976 (
            .O(N__23408),
            .I(N__23405));
    InMux I__2975 (
            .O(N__23405),
            .I(N__23402));
    LocalMux I__2974 (
            .O(N__23402),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__2973 (
            .O(N__23399),
            .I(N__23396));
    InMux I__2972 (
            .O(N__23396),
            .I(N__23393));
    LocalMux I__2971 (
            .O(N__23393),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__2970 (
            .O(N__23390),
            .I(N__23387));
    LocalMux I__2969 (
            .O(N__23387),
            .I(N__23384));
    Odrv4 I__2968 (
            .O(N__23384),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__2967 (
            .O(N__23381),
            .I(N__23378));
    InMux I__2966 (
            .O(N__23378),
            .I(N__23375));
    LocalMux I__2965 (
            .O(N__23375),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__2964 (
            .O(N__23372),
            .I(N__23369));
    LocalMux I__2963 (
            .O(N__23369),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__2962 (
            .O(N__23366),
            .I(N__23363));
    InMux I__2961 (
            .O(N__23363),
            .I(N__23360));
    LocalMux I__2960 (
            .O(N__23360),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__2959 (
            .O(N__23357),
            .I(N__23354));
    LocalMux I__2958 (
            .O(N__23354),
            .I(N__23351));
    Odrv4 I__2957 (
            .O(N__23351),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__2956 (
            .O(N__23348),
            .I(N__23345));
    InMux I__2955 (
            .O(N__23345),
            .I(N__23342));
    LocalMux I__2954 (
            .O(N__23342),
            .I(N__23339));
    Odrv4 I__2953 (
            .O(N__23339),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__2952 (
            .O(N__23336),
            .I(N__23333));
    LocalMux I__2951 (
            .O(N__23333),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__2950 (
            .O(N__23330),
            .I(N__23327));
    InMux I__2949 (
            .O(N__23327),
            .I(N__23324));
    LocalMux I__2948 (
            .O(N__23324),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__2947 (
            .O(N__23321),
            .I(N__23318));
    InMux I__2946 (
            .O(N__23318),
            .I(N__23315));
    LocalMux I__2945 (
            .O(N__23315),
            .I(N__23312));
    Odrv4 I__2944 (
            .O(N__23312),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__2943 (
            .O(N__23309),
            .I(N__23303));
    InMux I__2942 (
            .O(N__23308),
            .I(N__23303));
    LocalMux I__2941 (
            .O(N__23303),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__2940 (
            .O(N__23300),
            .I(N__23297));
    InMux I__2939 (
            .O(N__23297),
            .I(N__23291));
    InMux I__2938 (
            .O(N__23296),
            .I(N__23291));
    LocalMux I__2937 (
            .O(N__23291),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__2936 (
            .O(N__23288),
            .I(N__23284));
    InMux I__2935 (
            .O(N__23287),
            .I(N__23281));
    LocalMux I__2934 (
            .O(N__23284),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    LocalMux I__2933 (
            .O(N__23281),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2932 (
            .O(N__23276),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2931 (
            .O(N__23273),
            .I(N__23269));
    InMux I__2930 (
            .O(N__23272),
            .I(N__23266));
    LocalMux I__2929 (
            .O(N__23269),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    LocalMux I__2928 (
            .O(N__23266),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2927 (
            .O(N__23261),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2926 (
            .O(N__23258),
            .I(N__23255));
    LocalMux I__2925 (
            .O(N__23255),
            .I(N__23252));
    Span4Mux_h I__2924 (
            .O(N__23252),
            .I(N__23248));
    InMux I__2923 (
            .O(N__23251),
            .I(N__23245));
    Odrv4 I__2922 (
            .O(N__23248),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__2921 (
            .O(N__23245),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2920 (
            .O(N__23240),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    CascadeMux I__2919 (
            .O(N__23237),
            .I(N__23234));
    InMux I__2918 (
            .O(N__23234),
            .I(N__23230));
    InMux I__2917 (
            .O(N__23233),
            .I(N__23227));
    LocalMux I__2916 (
            .O(N__23230),
            .I(N__23222));
    LocalMux I__2915 (
            .O(N__23227),
            .I(N__23222));
    Odrv4 I__2914 (
            .O(N__23222),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2913 (
            .O(N__23219),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2912 (
            .O(N__23216),
            .I(N__23212));
    InMux I__2911 (
            .O(N__23215),
            .I(N__23209));
    LocalMux I__2910 (
            .O(N__23212),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    LocalMux I__2909 (
            .O(N__23209),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2908 (
            .O(N__23204),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2907 (
            .O(N__23201),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2906 (
            .O(N__23198),
            .I(N__23195));
    LocalMux I__2905 (
            .O(N__23195),
            .I(N__23192));
    Span4Mux_s2_h I__2904 (
            .O(N__23192),
            .I(N__23184));
    InMux I__2903 (
            .O(N__23191),
            .I(N__23179));
    InMux I__2902 (
            .O(N__23190),
            .I(N__23179));
    InMux I__2901 (
            .O(N__23189),
            .I(N__23176));
    InMux I__2900 (
            .O(N__23188),
            .I(N__23173));
    InMux I__2899 (
            .O(N__23187),
            .I(N__23170));
    Span4Mux_v I__2898 (
            .O(N__23184),
            .I(N__23155));
    LocalMux I__2897 (
            .O(N__23179),
            .I(N__23155));
    LocalMux I__2896 (
            .O(N__23176),
            .I(N__23155));
    LocalMux I__2895 (
            .O(N__23173),
            .I(N__23155));
    LocalMux I__2894 (
            .O(N__23170),
            .I(N__23155));
    InMux I__2893 (
            .O(N__23169),
            .I(N__23152));
    InMux I__2892 (
            .O(N__23168),
            .I(N__23147));
    InMux I__2891 (
            .O(N__23167),
            .I(N__23147));
    InMux I__2890 (
            .O(N__23166),
            .I(N__23144));
    Sp12to4 I__2889 (
            .O(N__23155),
            .I(N__23137));
    LocalMux I__2888 (
            .O(N__23152),
            .I(N__23137));
    LocalMux I__2887 (
            .O(N__23147),
            .I(N__23137));
    LocalMux I__2886 (
            .O(N__23144),
            .I(N__23134));
    Span12Mux_v I__2885 (
            .O(N__23137),
            .I(N__23131));
    Span12Mux_s5_h I__2884 (
            .O(N__23134),
            .I(N__23128));
    Odrv12 I__2883 (
            .O(N__23131),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv12 I__2882 (
            .O(N__23128),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__2881 (
            .O(N__23123),
            .I(N__23120));
    InMux I__2880 (
            .O(N__23120),
            .I(N__23117));
    LocalMux I__2879 (
            .O(N__23117),
            .I(N__23114));
    Odrv12 I__2878 (
            .O(N__23114),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__2877 (
            .O(N__23111),
            .I(N__23105));
    InMux I__2876 (
            .O(N__23110),
            .I(N__23105));
    LocalMux I__2875 (
            .O(N__23105),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2874 (
            .O(N__23102),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    CascadeMux I__2873 (
            .O(N__23099),
            .I(N__23096));
    InMux I__2872 (
            .O(N__23096),
            .I(N__23092));
    CascadeMux I__2871 (
            .O(N__23095),
            .I(N__23089));
    LocalMux I__2870 (
            .O(N__23092),
            .I(N__23086));
    InMux I__2869 (
            .O(N__23089),
            .I(N__23083));
    Odrv4 I__2868 (
            .O(N__23086),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    LocalMux I__2867 (
            .O(N__23083),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2866 (
            .O(N__23078),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    CascadeMux I__2865 (
            .O(N__23075),
            .I(N__23072));
    InMux I__2864 (
            .O(N__23072),
            .I(N__23068));
    InMux I__2863 (
            .O(N__23071),
            .I(N__23065));
    LocalMux I__2862 (
            .O(N__23068),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    LocalMux I__2861 (
            .O(N__23065),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2860 (
            .O(N__23060),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    CascadeMux I__2859 (
            .O(N__23057),
            .I(N__23053));
    InMux I__2858 (
            .O(N__23056),
            .I(N__23050));
    InMux I__2857 (
            .O(N__23053),
            .I(N__23047));
    LocalMux I__2856 (
            .O(N__23050),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    LocalMux I__2855 (
            .O(N__23047),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2854 (
            .O(N__23042),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__2853 (
            .O(N__23039),
            .I(N__23035));
    InMux I__2852 (
            .O(N__23038),
            .I(N__23032));
    LocalMux I__2851 (
            .O(N__23035),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__2850 (
            .O(N__23032),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2849 (
            .O(N__23027),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2848 (
            .O(N__23024),
            .I(N__23021));
    LocalMux I__2847 (
            .O(N__23021),
            .I(N__23017));
    InMux I__2846 (
            .O(N__23020),
            .I(N__23014));
    Odrv4 I__2845 (
            .O(N__23017),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    LocalMux I__2844 (
            .O(N__23014),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2843 (
            .O(N__23009),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2842 (
            .O(N__23006),
            .I(N__23000));
    InMux I__2841 (
            .O(N__23005),
            .I(N__23000));
    LocalMux I__2840 (
            .O(N__23000),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2839 (
            .O(N__22997),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    CascadeMux I__2838 (
            .O(N__22994),
            .I(N__22990));
    InMux I__2837 (
            .O(N__22993),
            .I(N__22985));
    InMux I__2836 (
            .O(N__22990),
            .I(N__22985));
    LocalMux I__2835 (
            .O(N__22985),
            .I(N__22982));
    Odrv4 I__2834 (
            .O(N__22982),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2833 (
            .O(N__22979),
            .I(bfn_5_18_0_));
    InMux I__2832 (
            .O(N__22976),
            .I(N__22972));
    InMux I__2831 (
            .O(N__22975),
            .I(N__22969));
    LocalMux I__2830 (
            .O(N__22972),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    LocalMux I__2829 (
            .O(N__22969),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2828 (
            .O(N__22964),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    InMux I__2827 (
            .O(N__22961),
            .I(N__22958));
    LocalMux I__2826 (
            .O(N__22958),
            .I(N__22953));
    InMux I__2825 (
            .O(N__22957),
            .I(N__22950));
    InMux I__2824 (
            .O(N__22956),
            .I(N__22947));
    Span4Mux_v I__2823 (
            .O(N__22953),
            .I(N__22940));
    LocalMux I__2822 (
            .O(N__22950),
            .I(N__22940));
    LocalMux I__2821 (
            .O(N__22947),
            .I(N__22940));
    Span4Mux_h I__2820 (
            .O(N__22940),
            .I(N__22937));
    Odrv4 I__2819 (
            .O(N__22937),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2818 (
            .O(N__22934),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    InMux I__2817 (
            .O(N__22931),
            .I(N__22928));
    LocalMux I__2816 (
            .O(N__22928),
            .I(N__22925));
    Odrv4 I__2815 (
            .O(N__22925),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__2814 (
            .O(N__22922),
            .I(N__22916));
    InMux I__2813 (
            .O(N__22921),
            .I(N__22916));
    LocalMux I__2812 (
            .O(N__22916),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2811 (
            .O(N__22913),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2810 (
            .O(N__22910),
            .I(N__22904));
    InMux I__2809 (
            .O(N__22909),
            .I(N__22904));
    LocalMux I__2808 (
            .O(N__22904),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2807 (
            .O(N__22901),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2806 (
            .O(N__22898),
            .I(N__22895));
    LocalMux I__2805 (
            .O(N__22895),
            .I(N__22892));
    Odrv12 I__2804 (
            .O(N__22892),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__2803 (
            .O(N__22889),
            .I(N__22886));
    LocalMux I__2802 (
            .O(N__22886),
            .I(N__22882));
    InMux I__2801 (
            .O(N__22885),
            .I(N__22879));
    Odrv4 I__2800 (
            .O(N__22882),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    LocalMux I__2799 (
            .O(N__22879),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2798 (
            .O(N__22874),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2797 (
            .O(N__22871),
            .I(N__22868));
    LocalMux I__2796 (
            .O(N__22868),
            .I(N__22865));
    Odrv4 I__2795 (
            .O(N__22865),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    InMux I__2794 (
            .O(N__22862),
            .I(N__22856));
    InMux I__2793 (
            .O(N__22861),
            .I(N__22856));
    LocalMux I__2792 (
            .O(N__22856),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2791 (
            .O(N__22853),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2790 (
            .O(N__22850),
            .I(N__22846));
    InMux I__2789 (
            .O(N__22849),
            .I(N__22843));
    LocalMux I__2788 (
            .O(N__22846),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    LocalMux I__2787 (
            .O(N__22843),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2786 (
            .O(N__22838),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2785 (
            .O(N__22835),
            .I(N__22831));
    InMux I__2784 (
            .O(N__22834),
            .I(N__22828));
    LocalMux I__2783 (
            .O(N__22831),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2782 (
            .O(N__22828),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2781 (
            .O(N__22823),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    CascadeMux I__2780 (
            .O(N__22820),
            .I(N__22817));
    InMux I__2779 (
            .O(N__22817),
            .I(N__22813));
    InMux I__2778 (
            .O(N__22816),
            .I(N__22810));
    LocalMux I__2777 (
            .O(N__22813),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    LocalMux I__2776 (
            .O(N__22810),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2775 (
            .O(N__22805),
            .I(bfn_5_17_0_));
    InMux I__2774 (
            .O(N__22802),
            .I(N__22799));
    LocalMux I__2773 (
            .O(N__22799),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__2772 (
            .O(N__22796),
            .I(N__22793));
    LocalMux I__2771 (
            .O(N__22793),
            .I(N__22790));
    Span4Mux_h I__2770 (
            .O(N__22790),
            .I(N__22787));
    Odrv4 I__2769 (
            .O(N__22787),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2768 (
            .O(N__22784),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    InMux I__2767 (
            .O(N__22781),
            .I(N__22778));
    LocalMux I__2766 (
            .O(N__22778),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__2765 (
            .O(N__22775),
            .I(N__22772));
    LocalMux I__2764 (
            .O(N__22772),
            .I(N__22769));
    Span4Mux_h I__2763 (
            .O(N__22769),
            .I(N__22766));
    Odrv4 I__2762 (
            .O(N__22766),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2761 (
            .O(N__22763),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    CascadeMux I__2760 (
            .O(N__22760),
            .I(N__22757));
    InMux I__2759 (
            .O(N__22757),
            .I(N__22754));
    LocalMux I__2758 (
            .O(N__22754),
            .I(N__22749));
    InMux I__2757 (
            .O(N__22753),
            .I(N__22746));
    InMux I__2756 (
            .O(N__22752),
            .I(N__22743));
    Span4Mux_v I__2755 (
            .O(N__22749),
            .I(N__22738));
    LocalMux I__2754 (
            .O(N__22746),
            .I(N__22738));
    LocalMux I__2753 (
            .O(N__22743),
            .I(N__22735));
    Span4Mux_h I__2752 (
            .O(N__22738),
            .I(N__22732));
    Span4Mux_h I__2751 (
            .O(N__22735),
            .I(N__22729));
    Odrv4 I__2750 (
            .O(N__22732),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__2749 (
            .O(N__22729),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2748 (
            .O(N__22724),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    CascadeMux I__2747 (
            .O(N__22721),
            .I(N__22718));
    InMux I__2746 (
            .O(N__22718),
            .I(N__22715));
    LocalMux I__2745 (
            .O(N__22715),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__2744 (
            .O(N__22712),
            .I(N__22708));
    InMux I__2743 (
            .O(N__22711),
            .I(N__22704));
    InMux I__2742 (
            .O(N__22708),
            .I(N__22698));
    InMux I__2741 (
            .O(N__22707),
            .I(N__22698));
    LocalMux I__2740 (
            .O(N__22704),
            .I(N__22695));
    InMux I__2739 (
            .O(N__22703),
            .I(N__22692));
    LocalMux I__2738 (
            .O(N__22698),
            .I(N__22689));
    Span4Mux_h I__2737 (
            .O(N__22695),
            .I(N__22686));
    LocalMux I__2736 (
            .O(N__22692),
            .I(N__22683));
    Span4Mux_v I__2735 (
            .O(N__22689),
            .I(N__22680));
    Span4Mux_v I__2734 (
            .O(N__22686),
            .I(N__22675));
    Span4Mux_h I__2733 (
            .O(N__22683),
            .I(N__22675));
    Odrv4 I__2732 (
            .O(N__22680),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2731 (
            .O(N__22675),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2730 (
            .O(N__22670),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2729 (
            .O(N__22667),
            .I(N__22664));
    LocalMux I__2728 (
            .O(N__22664),
            .I(N__22661));
    Odrv4 I__2727 (
            .O(N__22661),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__2726 (
            .O(N__22658),
            .I(N__22655));
    LocalMux I__2725 (
            .O(N__22655),
            .I(N__22651));
    InMux I__2724 (
            .O(N__22654),
            .I(N__22648));
    Span4Mux_v I__2723 (
            .O(N__22651),
            .I(N__22642));
    LocalMux I__2722 (
            .O(N__22648),
            .I(N__22642));
    InMux I__2721 (
            .O(N__22647),
            .I(N__22639));
    Span4Mux_h I__2720 (
            .O(N__22642),
            .I(N__22636));
    LocalMux I__2719 (
            .O(N__22639),
            .I(N__22633));
    Odrv4 I__2718 (
            .O(N__22636),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__2717 (
            .O(N__22633),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2716 (
            .O(N__22628),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2715 (
            .O(N__22625),
            .I(N__22622));
    LocalMux I__2714 (
            .O(N__22622),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__2713 (
            .O(N__22619),
            .I(N__22616));
    InMux I__2712 (
            .O(N__22616),
            .I(N__22613));
    LocalMux I__2711 (
            .O(N__22613),
            .I(N__22609));
    InMux I__2710 (
            .O(N__22612),
            .I(N__22606));
    Span4Mux_h I__2709 (
            .O(N__22609),
            .I(N__22602));
    LocalMux I__2708 (
            .O(N__22606),
            .I(N__22599));
    InMux I__2707 (
            .O(N__22605),
            .I(N__22596));
    Span4Mux_v I__2706 (
            .O(N__22602),
            .I(N__22593));
    Span4Mux_h I__2705 (
            .O(N__22599),
            .I(N__22590));
    LocalMux I__2704 (
            .O(N__22596),
            .I(N__22587));
    Odrv4 I__2703 (
            .O(N__22593),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2702 (
            .O(N__22590),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2701 (
            .O(N__22587),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2700 (
            .O(N__22580),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__2699 (
            .O(N__22577),
            .I(N__22574));
    LocalMux I__2698 (
            .O(N__22574),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__2697 (
            .O(N__22571),
            .I(N__22568));
    InMux I__2696 (
            .O(N__22568),
            .I(N__22565));
    LocalMux I__2695 (
            .O(N__22565),
            .I(N__22560));
    InMux I__2694 (
            .O(N__22564),
            .I(N__22557));
    InMux I__2693 (
            .O(N__22563),
            .I(N__22554));
    Span4Mux_v I__2692 (
            .O(N__22560),
            .I(N__22547));
    LocalMux I__2691 (
            .O(N__22557),
            .I(N__22547));
    LocalMux I__2690 (
            .O(N__22554),
            .I(N__22547));
    Span4Mux_h I__2689 (
            .O(N__22547),
            .I(N__22544));
    Odrv4 I__2688 (
            .O(N__22544),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2687 (
            .O(N__22541),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2686 (
            .O(N__22538),
            .I(N__22534));
    InMux I__2685 (
            .O(N__22537),
            .I(N__22531));
    LocalMux I__2684 (
            .O(N__22534),
            .I(N__22527));
    LocalMux I__2683 (
            .O(N__22531),
            .I(N__22524));
    InMux I__2682 (
            .O(N__22530),
            .I(N__22521));
    Span4Mux_h I__2681 (
            .O(N__22527),
            .I(N__22518));
    Span4Mux_h I__2680 (
            .O(N__22524),
            .I(N__22513));
    LocalMux I__2679 (
            .O(N__22521),
            .I(N__22513));
    Odrv4 I__2678 (
            .O(N__22518),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2677 (
            .O(N__22513),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2676 (
            .O(N__22508),
            .I(bfn_5_16_0_));
    InMux I__2675 (
            .O(N__22505),
            .I(N__22502));
    LocalMux I__2674 (
            .O(N__22502),
            .I(N__22499));
    Span4Mux_h I__2673 (
            .O(N__22499),
            .I(N__22496));
    Odrv4 I__2672 (
            .O(N__22496),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2671 (
            .O(N__22493),
            .I(N__22490));
    LocalMux I__2670 (
            .O(N__22490),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ));
    InMux I__2669 (
            .O(N__22487),
            .I(N__22484));
    LocalMux I__2668 (
            .O(N__22484),
            .I(N__22481));
    Odrv12 I__2667 (
            .O(N__22481),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    CascadeMux I__2666 (
            .O(N__22478),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_ ));
    InMux I__2665 (
            .O(N__22475),
            .I(N__22471));
    InMux I__2664 (
            .O(N__22474),
            .I(N__22468));
    LocalMux I__2663 (
            .O(N__22471),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    LocalMux I__2662 (
            .O(N__22468),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    InMux I__2661 (
            .O(N__22463),
            .I(N__22457));
    InMux I__2660 (
            .O(N__22462),
            .I(N__22457));
    LocalMux I__2659 (
            .O(N__22457),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    InMux I__2658 (
            .O(N__22454),
            .I(N__22451));
    LocalMux I__2657 (
            .O(N__22451),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    CascadeMux I__2656 (
            .O(N__22448),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ));
    InMux I__2655 (
            .O(N__22445),
            .I(N__22442));
    LocalMux I__2654 (
            .O(N__22442),
            .I(N__22439));
    Odrv4 I__2653 (
            .O(N__22439),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    CascadeMux I__2652 (
            .O(N__22436),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ));
    CascadeMux I__2651 (
            .O(N__22433),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ));
    InMux I__2650 (
            .O(N__22430),
            .I(N__22427));
    LocalMux I__2649 (
            .O(N__22427),
            .I(N__22424));
    Odrv12 I__2648 (
            .O(N__22424),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    CascadeMux I__2647 (
            .O(N__22421),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ));
    InMux I__2646 (
            .O(N__22418),
            .I(N__22415));
    LocalMux I__2645 (
            .O(N__22415),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    CascadeMux I__2644 (
            .O(N__22412),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ));
    InMux I__2643 (
            .O(N__22409),
            .I(N__22401));
    CascadeMux I__2642 (
            .O(N__22408),
            .I(N__22398));
    InMux I__2641 (
            .O(N__22407),
            .I(N__22395));
    InMux I__2640 (
            .O(N__22406),
            .I(N__22388));
    InMux I__2639 (
            .O(N__22405),
            .I(N__22388));
    InMux I__2638 (
            .O(N__22404),
            .I(N__22388));
    LocalMux I__2637 (
            .O(N__22401),
            .I(N__22385));
    InMux I__2636 (
            .O(N__22398),
            .I(N__22382));
    LocalMux I__2635 (
            .O(N__22395),
            .I(N__22377));
    LocalMux I__2634 (
            .O(N__22388),
            .I(N__22377));
    Span4Mux_v I__2633 (
            .O(N__22385),
            .I(N__22373));
    LocalMux I__2632 (
            .O(N__22382),
            .I(N__22368));
    Span4Mux_v I__2631 (
            .O(N__22377),
            .I(N__22368));
    InMux I__2630 (
            .O(N__22376),
            .I(N__22365));
    Span4Mux_v I__2629 (
            .O(N__22373),
            .I(N__22362));
    Span4Mux_h I__2628 (
            .O(N__22368),
            .I(N__22359));
    LocalMux I__2627 (
            .O(N__22365),
            .I(N__22356));
    Odrv4 I__2626 (
            .O(N__22362),
            .I(\current_shift_inst.PI_CTRL.N_164 ));
    Odrv4 I__2625 (
            .O(N__22359),
            .I(\current_shift_inst.PI_CTRL.N_164 ));
    Odrv4 I__2624 (
            .O(N__22356),
            .I(\current_shift_inst.PI_CTRL.N_164 ));
    InMux I__2623 (
            .O(N__22349),
            .I(N__22346));
    LocalMux I__2622 (
            .O(N__22346),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    CascadeMux I__2621 (
            .O(N__22343),
            .I(N__22340));
    InMux I__2620 (
            .O(N__22340),
            .I(N__22337));
    LocalMux I__2619 (
            .O(N__22337),
            .I(N__22334));
    Odrv4 I__2618 (
            .O(N__22334),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__2617 (
            .O(N__22331),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ));
    InMux I__2616 (
            .O(N__22328),
            .I(N__22325));
    LocalMux I__2615 (
            .O(N__22325),
            .I(N__22322));
    Odrv4 I__2614 (
            .O(N__22322),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    CascadeMux I__2613 (
            .O(N__22319),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    InMux I__2612 (
            .O(N__22316),
            .I(N__22313));
    LocalMux I__2611 (
            .O(N__22313),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__2610 (
            .O(N__22310),
            .I(N__22307));
    LocalMux I__2609 (
            .O(N__22307),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__2608 (
            .O(N__22304),
            .I(N__22300));
    CascadeMux I__2607 (
            .O(N__22303),
            .I(N__22297));
    InMux I__2606 (
            .O(N__22300),
            .I(N__22288));
    InMux I__2605 (
            .O(N__22297),
            .I(N__22288));
    InMux I__2604 (
            .O(N__22296),
            .I(N__22285));
    InMux I__2603 (
            .O(N__22295),
            .I(N__22282));
    InMux I__2602 (
            .O(N__22294),
            .I(N__22276));
    InMux I__2601 (
            .O(N__22293),
            .I(N__22273));
    LocalMux I__2600 (
            .O(N__22288),
            .I(N__22266));
    LocalMux I__2599 (
            .O(N__22285),
            .I(N__22266));
    LocalMux I__2598 (
            .O(N__22282),
            .I(N__22266));
    InMux I__2597 (
            .O(N__22281),
            .I(N__22261));
    InMux I__2596 (
            .O(N__22280),
            .I(N__22261));
    InMux I__2595 (
            .O(N__22279),
            .I(N__22258));
    LocalMux I__2594 (
            .O(N__22276),
            .I(N__22253));
    LocalMux I__2593 (
            .O(N__22273),
            .I(N__22253));
    Span4Mux_s3_h I__2592 (
            .O(N__22266),
            .I(N__22250));
    LocalMux I__2591 (
            .O(N__22261),
            .I(N__22247));
    LocalMux I__2590 (
            .O(N__22258),
            .I(N__22244));
    Span4Mux_v I__2589 (
            .O(N__22253),
            .I(N__22241));
    Span4Mux_v I__2588 (
            .O(N__22250),
            .I(N__22236));
    Span4Mux_v I__2587 (
            .O(N__22247),
            .I(N__22236));
    Span4Mux_h I__2586 (
            .O(N__22244),
            .I(N__22233));
    Odrv4 I__2585 (
            .O(N__22241),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2584 (
            .O(N__22236),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2583 (
            .O(N__22233),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    InMux I__2582 (
            .O(N__22226),
            .I(N__22223));
    LocalMux I__2581 (
            .O(N__22223),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    CascadeMux I__2580 (
            .O(N__22220),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ));
    InMux I__2579 (
            .O(N__22217),
            .I(N__22214));
    LocalMux I__2578 (
            .O(N__22214),
            .I(\current_shift_inst.PI_CTRL.N_71 ));
    CascadeMux I__2577 (
            .O(N__22211),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ));
    InMux I__2576 (
            .O(N__22208),
            .I(N__22205));
    LocalMux I__2575 (
            .O(N__22205),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ));
    InMux I__2574 (
            .O(N__22202),
            .I(N__22199));
    LocalMux I__2573 (
            .O(N__22199),
            .I(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ));
    IoInMux I__2572 (
            .O(N__22196),
            .I(N__22193));
    LocalMux I__2571 (
            .O(N__22193),
            .I(N__22190));
    Span4Mux_s1_v I__2570 (
            .O(N__22190),
            .I(N__22187));
    Sp12to4 I__2569 (
            .O(N__22187),
            .I(N__22184));
    Span12Mux_s10_h I__2568 (
            .O(N__22184),
            .I(N__22181));
    Span12Mux_h I__2567 (
            .O(N__22181),
            .I(N__22178));
    Span12Mux_v I__2566 (
            .O(N__22178),
            .I(N__22175));
    Odrv12 I__2565 (
            .O(N__22175),
            .I(pwm_output_c));
    CascadeMux I__2564 (
            .O(N__22172),
            .I(N__22169));
    InMux I__2563 (
            .O(N__22169),
            .I(N__22166));
    LocalMux I__2562 (
            .O(N__22166),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671 ));
    CascadeMux I__2561 (
            .O(N__22163),
            .I(N__22160));
    InMux I__2560 (
            .O(N__22160),
            .I(N__22157));
    LocalMux I__2559 (
            .O(N__22157),
            .I(\pwm_generator_inst.threshold_9 ));
    CascadeMux I__2558 (
            .O(N__22154),
            .I(N__22151));
    InMux I__2557 (
            .O(N__22151),
            .I(N__22148));
    LocalMux I__2556 (
            .O(N__22148),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271 ));
    CascadeMux I__2555 (
            .O(N__22145),
            .I(N__22142));
    InMux I__2554 (
            .O(N__22142),
            .I(N__22139));
    LocalMux I__2553 (
            .O(N__22139),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__2552 (
            .O(N__22136),
            .I(N__22133));
    LocalMux I__2551 (
            .O(N__22133),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61 ));
    CascadeMux I__2550 (
            .O(N__22130),
            .I(N__22127));
    InMux I__2549 (
            .O(N__22127),
            .I(N__22124));
    LocalMux I__2548 (
            .O(N__22124),
            .I(N__22121));
    Odrv4 I__2547 (
            .O(N__22121),
            .I(\pwm_generator_inst.un14_counter_7 ));
    CascadeMux I__2546 (
            .O(N__22118),
            .I(N__22111));
    InMux I__2545 (
            .O(N__22117),
            .I(N__22100));
    InMux I__2544 (
            .O(N__22116),
            .I(N__22100));
    InMux I__2543 (
            .O(N__22115),
            .I(N__22100));
    InMux I__2542 (
            .O(N__22114),
            .I(N__22100));
    InMux I__2541 (
            .O(N__22111),
            .I(N__22094));
    InMux I__2540 (
            .O(N__22110),
            .I(N__22089));
    InMux I__2539 (
            .O(N__22109),
            .I(N__22089));
    LocalMux I__2538 (
            .O(N__22100),
            .I(N__22086));
    InMux I__2537 (
            .O(N__22099),
            .I(N__22079));
    InMux I__2536 (
            .O(N__22098),
            .I(N__22079));
    InMux I__2535 (
            .O(N__22097),
            .I(N__22079));
    LocalMux I__2534 (
            .O(N__22094),
            .I(N__22074));
    LocalMux I__2533 (
            .O(N__22089),
            .I(N__22074));
    Span4Mux_v I__2532 (
            .O(N__22086),
            .I(N__22069));
    LocalMux I__2531 (
            .O(N__22079),
            .I(N__22069));
    Span4Mux_v I__2530 (
            .O(N__22074),
            .I(N__22066));
    Odrv4 I__2529 (
            .O(N__22069),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2528 (
            .O(N__22066),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__2527 (
            .O(N__22061),
            .I(N__22054));
    CascadeMux I__2526 (
            .O(N__22060),
            .I(N__22050));
    CascadeMux I__2525 (
            .O(N__22059),
            .I(N__22045));
    CascadeMux I__2524 (
            .O(N__22058),
            .I(N__22041));
    CascadeMux I__2523 (
            .O(N__22057),
            .I(N__22037));
    InMux I__2522 (
            .O(N__22054),
            .I(N__22032));
    InMux I__2521 (
            .O(N__22053),
            .I(N__22032));
    InMux I__2520 (
            .O(N__22050),
            .I(N__22029));
    InMux I__2519 (
            .O(N__22049),
            .I(N__22020));
    InMux I__2518 (
            .O(N__22048),
            .I(N__22020));
    InMux I__2517 (
            .O(N__22045),
            .I(N__22020));
    InMux I__2516 (
            .O(N__22044),
            .I(N__22020));
    InMux I__2515 (
            .O(N__22041),
            .I(N__22013));
    InMux I__2514 (
            .O(N__22040),
            .I(N__22013));
    InMux I__2513 (
            .O(N__22037),
            .I(N__22013));
    LocalMux I__2512 (
            .O(N__22032),
            .I(N__21999));
    LocalMux I__2511 (
            .O(N__22029),
            .I(N__21999));
    LocalMux I__2510 (
            .O(N__22020),
            .I(N__21999));
    LocalMux I__2509 (
            .O(N__22013),
            .I(N__21999));
    InMux I__2508 (
            .O(N__22012),
            .I(N__21979));
    InMux I__2507 (
            .O(N__22011),
            .I(N__21979));
    InMux I__2506 (
            .O(N__22010),
            .I(N__21972));
    InMux I__2505 (
            .O(N__22009),
            .I(N__21972));
    InMux I__2504 (
            .O(N__22008),
            .I(N__21972));
    Span4Mux_v I__2503 (
            .O(N__21999),
            .I(N__21969));
    InMux I__2502 (
            .O(N__21998),
            .I(N__21951));
    InMux I__2501 (
            .O(N__21997),
            .I(N__21951));
    InMux I__2500 (
            .O(N__21996),
            .I(N__21951));
    InMux I__2499 (
            .O(N__21995),
            .I(N__21951));
    InMux I__2498 (
            .O(N__21994),
            .I(N__21951));
    InMux I__2497 (
            .O(N__21993),
            .I(N__21951));
    InMux I__2496 (
            .O(N__21992),
            .I(N__21951));
    InMux I__2495 (
            .O(N__21991),
            .I(N__21951));
    InMux I__2494 (
            .O(N__21990),
            .I(N__21936));
    InMux I__2493 (
            .O(N__21989),
            .I(N__21936));
    InMux I__2492 (
            .O(N__21988),
            .I(N__21936));
    InMux I__2491 (
            .O(N__21987),
            .I(N__21936));
    InMux I__2490 (
            .O(N__21986),
            .I(N__21936));
    InMux I__2489 (
            .O(N__21985),
            .I(N__21936));
    InMux I__2488 (
            .O(N__21984),
            .I(N__21936));
    LocalMux I__2487 (
            .O(N__21979),
            .I(N__21931));
    LocalMux I__2486 (
            .O(N__21972),
            .I(N__21931));
    Span4Mux_v I__2485 (
            .O(N__21969),
            .I(N__21928));
    CascadeMux I__2484 (
            .O(N__21968),
            .I(N__21925));
    LocalMux I__2483 (
            .O(N__21951),
            .I(N__21917));
    LocalMux I__2482 (
            .O(N__21936),
            .I(N__21917));
    Span4Mux_v I__2481 (
            .O(N__21931),
            .I(N__21917));
    Span4Mux_v I__2480 (
            .O(N__21928),
            .I(N__21914));
    InMux I__2479 (
            .O(N__21925),
            .I(N__21911));
    InMux I__2478 (
            .O(N__21924),
            .I(N__21908));
    Span4Mux_v I__2477 (
            .O(N__21917),
            .I(N__21905));
    Odrv4 I__2476 (
            .O(N__21914),
            .I(N_19_1));
    LocalMux I__2475 (
            .O(N__21911),
            .I(N_19_1));
    LocalMux I__2474 (
            .O(N__21908),
            .I(N_19_1));
    Odrv4 I__2473 (
            .O(N__21905),
            .I(N_19_1));
    CascadeMux I__2472 (
            .O(N__21896),
            .I(N__21893));
    InMux I__2471 (
            .O(N__21893),
            .I(N__21890));
    LocalMux I__2470 (
            .O(N__21890),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1 ));
    InMux I__2469 (
            .O(N__21887),
            .I(N__21872));
    InMux I__2468 (
            .O(N__21886),
            .I(N__21872));
    InMux I__2467 (
            .O(N__21885),
            .I(N__21872));
    InMux I__2466 (
            .O(N__21884),
            .I(N__21872));
    InMux I__2465 (
            .O(N__21883),
            .I(N__21865));
    InMux I__2464 (
            .O(N__21882),
            .I(N__21865));
    InMux I__2463 (
            .O(N__21881),
            .I(N__21865));
    LocalMux I__2462 (
            .O(N__21872),
            .I(N__21857));
    LocalMux I__2461 (
            .O(N__21865),
            .I(N__21857));
    InMux I__2460 (
            .O(N__21864),
            .I(N__21850));
    InMux I__2459 (
            .O(N__21863),
            .I(N__21850));
    InMux I__2458 (
            .O(N__21862),
            .I(N__21850));
    Span4Mux_v I__2457 (
            .O(N__21857),
            .I(N__21845));
    LocalMux I__2456 (
            .O(N__21850),
            .I(N__21845));
    Span4Mux_v I__2455 (
            .O(N__21845),
            .I(N__21842));
    Odrv4 I__2454 (
            .O(N__21842),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__2453 (
            .O(N__21839),
            .I(N__21836));
    InMux I__2452 (
            .O(N__21836),
            .I(N__21833));
    LocalMux I__2451 (
            .O(N__21833),
            .I(N__21830));
    Odrv4 I__2450 (
            .O(N__21830),
            .I(\pwm_generator_inst.threshold_3 ));
    CascadeMux I__2449 (
            .O(N__21827),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ));
    CascadeMux I__2448 (
            .O(N__21824),
            .I(N__21821));
    InMux I__2447 (
            .O(N__21821),
            .I(N__21818));
    LocalMux I__2446 (
            .O(N__21818),
            .I(N__21815));
    Span4Mux_v I__2445 (
            .O(N__21815),
            .I(N__21811));
    InMux I__2444 (
            .O(N__21814),
            .I(N__21808));
    Odrv4 I__2443 (
            .O(N__21811),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__2442 (
            .O(N__21808),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__2441 (
            .O(N__21803),
            .I(N__21800));
    LocalMux I__2440 (
            .O(N__21800),
            .I(N__21796));
    InMux I__2439 (
            .O(N__21799),
            .I(N__21792));
    Span4Mux_v I__2438 (
            .O(N__21796),
            .I(N__21789));
    InMux I__2437 (
            .O(N__21795),
            .I(N__21786));
    LocalMux I__2436 (
            .O(N__21792),
            .I(N__21781));
    Span4Mux_v I__2435 (
            .O(N__21789),
            .I(N__21781));
    LocalMux I__2434 (
            .O(N__21786),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__2433 (
            .O(N__21781),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__2432 (
            .O(N__21776),
            .I(N__21773));
    LocalMux I__2431 (
            .O(N__21773),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__2430 (
            .O(N__21770),
            .I(N__21767));
    InMux I__2429 (
            .O(N__21767),
            .I(N__21764));
    LocalMux I__2428 (
            .O(N__21764),
            .I(\pwm_generator_inst.threshold_4 ));
    InMux I__2427 (
            .O(N__21761),
            .I(N__21758));
    LocalMux I__2426 (
            .O(N__21758),
            .I(N__21754));
    InMux I__2425 (
            .O(N__21757),
            .I(N__21750));
    Span4Mux_h I__2424 (
            .O(N__21754),
            .I(N__21747));
    InMux I__2423 (
            .O(N__21753),
            .I(N__21744));
    LocalMux I__2422 (
            .O(N__21750),
            .I(N__21741));
    Span4Mux_v I__2421 (
            .O(N__21747),
            .I(N__21738));
    LocalMux I__2420 (
            .O(N__21744),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv12 I__2419 (
            .O(N__21741),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__2418 (
            .O(N__21738),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__2417 (
            .O(N__21731),
            .I(N__21728));
    LocalMux I__2416 (
            .O(N__21728),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__2415 (
            .O(N__21725),
            .I(N__21722));
    InMux I__2414 (
            .O(N__21722),
            .I(N__21719));
    LocalMux I__2413 (
            .O(N__21719),
            .I(\pwm_generator_inst.threshold_5 ));
    InMux I__2412 (
            .O(N__21716),
            .I(N__21712));
    InMux I__2411 (
            .O(N__21715),
            .I(N__21709));
    LocalMux I__2410 (
            .O(N__21712),
            .I(N__21706));
    LocalMux I__2409 (
            .O(N__21709),
            .I(N__21703));
    Span4Mux_h I__2408 (
            .O(N__21706),
            .I(N__21699));
    Span4Mux_v I__2407 (
            .O(N__21703),
            .I(N__21696));
    InMux I__2406 (
            .O(N__21702),
            .I(N__21693));
    Span4Mux_v I__2405 (
            .O(N__21699),
            .I(N__21690));
    Odrv4 I__2404 (
            .O(N__21696),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2403 (
            .O(N__21693),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__2402 (
            .O(N__21690),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2401 (
            .O(N__21683),
            .I(N__21680));
    LocalMux I__2400 (
            .O(N__21680),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__2399 (
            .O(N__21677),
            .I(N__21674));
    InMux I__2398 (
            .O(N__21674),
            .I(N__21671));
    LocalMux I__2397 (
            .O(N__21671),
            .I(N__21668));
    Odrv4 I__2396 (
            .O(N__21668),
            .I(\pwm_generator_inst.un14_counter_6 ));
    InMux I__2395 (
            .O(N__21665),
            .I(N__21661));
    InMux I__2394 (
            .O(N__21664),
            .I(N__21658));
    LocalMux I__2393 (
            .O(N__21661),
            .I(N__21655));
    LocalMux I__2392 (
            .O(N__21658),
            .I(N__21651));
    Span4Mux_h I__2391 (
            .O(N__21655),
            .I(N__21648));
    InMux I__2390 (
            .O(N__21654),
            .I(N__21645));
    Span12Mux_h I__2389 (
            .O(N__21651),
            .I(N__21642));
    Odrv4 I__2388 (
            .O(N__21648),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2387 (
            .O(N__21645),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv12 I__2386 (
            .O(N__21642),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__2385 (
            .O(N__21635),
            .I(N__21632));
    LocalMux I__2384 (
            .O(N__21632),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__2383 (
            .O(N__21629),
            .I(N__21625));
    InMux I__2382 (
            .O(N__21628),
            .I(N__21622));
    LocalMux I__2381 (
            .O(N__21625),
            .I(N__21619));
    LocalMux I__2380 (
            .O(N__21622),
            .I(N__21615));
    Span4Mux_h I__2379 (
            .O(N__21619),
            .I(N__21612));
    InMux I__2378 (
            .O(N__21618),
            .I(N__21609));
    Span4Mux_h I__2377 (
            .O(N__21615),
            .I(N__21606));
    Span4Mux_v I__2376 (
            .O(N__21612),
            .I(N__21603));
    LocalMux I__2375 (
            .O(N__21609),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2374 (
            .O(N__21606),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2373 (
            .O(N__21603),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__2372 (
            .O(N__21596),
            .I(N__21593));
    LocalMux I__2371 (
            .O(N__21593),
            .I(\pwm_generator_inst.counter_i_7 ));
    InMux I__2370 (
            .O(N__21590),
            .I(N__21587));
    LocalMux I__2369 (
            .O(N__21587),
            .I(N__21583));
    InMux I__2368 (
            .O(N__21586),
            .I(N__21579));
    Span4Mux_v I__2367 (
            .O(N__21583),
            .I(N__21576));
    InMux I__2366 (
            .O(N__21582),
            .I(N__21573));
    LocalMux I__2365 (
            .O(N__21579),
            .I(N__21566));
    Span4Mux_v I__2364 (
            .O(N__21576),
            .I(N__21566));
    LocalMux I__2363 (
            .O(N__21573),
            .I(N__21566));
    Odrv4 I__2362 (
            .O(N__21566),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2361 (
            .O(N__21563),
            .I(N__21560));
    LocalMux I__2360 (
            .O(N__21560),
            .I(\pwm_generator_inst.counter_i_8 ));
    InMux I__2359 (
            .O(N__21557),
            .I(N__21554));
    LocalMux I__2358 (
            .O(N__21554),
            .I(N__21551));
    Span4Mux_v I__2357 (
            .O(N__21551),
            .I(N__21546));
    InMux I__2356 (
            .O(N__21550),
            .I(N__21543));
    InMux I__2355 (
            .O(N__21549),
            .I(N__21540));
    Span4Mux_v I__2354 (
            .O(N__21546),
            .I(N__21535));
    LocalMux I__2353 (
            .O(N__21543),
            .I(N__21535));
    LocalMux I__2352 (
            .O(N__21540),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__2351 (
            .O(N__21535),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__2350 (
            .O(N__21530),
            .I(N__21527));
    LocalMux I__2349 (
            .O(N__21527),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2348 (
            .O(N__21524),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    InMux I__2347 (
            .O(N__21521),
            .I(N__21503));
    InMux I__2346 (
            .O(N__21520),
            .I(N__21503));
    InMux I__2345 (
            .O(N__21519),
            .I(N__21503));
    InMux I__2344 (
            .O(N__21518),
            .I(N__21503));
    InMux I__2343 (
            .O(N__21517),
            .I(N__21494));
    InMux I__2342 (
            .O(N__21516),
            .I(N__21494));
    InMux I__2341 (
            .O(N__21515),
            .I(N__21494));
    InMux I__2340 (
            .O(N__21514),
            .I(N__21494));
    InMux I__2339 (
            .O(N__21513),
            .I(N__21489));
    InMux I__2338 (
            .O(N__21512),
            .I(N__21489));
    LocalMux I__2337 (
            .O(N__21503),
            .I(N__21484));
    LocalMux I__2336 (
            .O(N__21494),
            .I(N__21484));
    LocalMux I__2335 (
            .O(N__21489),
            .I(N__21481));
    Span4Mux_s3_h I__2334 (
            .O(N__21484),
            .I(N__21478));
    Odrv4 I__2333 (
            .O(N__21481),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__2332 (
            .O(N__21478),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__2331 (
            .O(N__21473),
            .I(N__21467));
    InMux I__2330 (
            .O(N__21472),
            .I(N__21460));
    InMux I__2329 (
            .O(N__21471),
            .I(N__21460));
    InMux I__2328 (
            .O(N__21470),
            .I(N__21460));
    LocalMux I__2327 (
            .O(N__21467),
            .I(N__21457));
    LocalMux I__2326 (
            .O(N__21460),
            .I(N__21454));
    Span4Mux_s3_h I__2325 (
            .O(N__21457),
            .I(N__21450));
    Span4Mux_s3_h I__2324 (
            .O(N__21454),
            .I(N__21447));
    InMux I__2323 (
            .O(N__21453),
            .I(N__21444));
    Odrv4 I__2322 (
            .O(N__21450),
            .I(\current_shift_inst.PI_CTRL.N_144 ));
    Odrv4 I__2321 (
            .O(N__21447),
            .I(\current_shift_inst.PI_CTRL.N_144 ));
    LocalMux I__2320 (
            .O(N__21444),
            .I(\current_shift_inst.PI_CTRL.N_144 ));
    InMux I__2319 (
            .O(N__21437),
            .I(N__21434));
    LocalMux I__2318 (
            .O(N__21434),
            .I(N__21431));
    Odrv4 I__2317 (
            .O(N__21431),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1 ));
    InMux I__2316 (
            .O(N__21428),
            .I(N__21425));
    LocalMux I__2315 (
            .O(N__21425),
            .I(N__21422));
    Odrv4 I__2314 (
            .O(N__21422),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31 ));
    CascadeMux I__2313 (
            .O(N__21419),
            .I(N__21416));
    InMux I__2312 (
            .O(N__21416),
            .I(N__21413));
    LocalMux I__2311 (
            .O(N__21413),
            .I(\current_shift_inst.PI_CTRL.N_146 ));
    CascadeMux I__2310 (
            .O(N__21410),
            .I(N__21407));
    InMux I__2309 (
            .O(N__21407),
            .I(N__21404));
    LocalMux I__2308 (
            .O(N__21404),
            .I(N__21401));
    Span4Mux_h I__2307 (
            .O(N__21401),
            .I(N__21398));
    Odrv4 I__2306 (
            .O(N__21398),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61 ));
    CascadeMux I__2305 (
            .O(N__21395),
            .I(N__21392));
    InMux I__2304 (
            .O(N__21392),
            .I(N__21389));
    LocalMux I__2303 (
            .O(N__21389),
            .I(N__21386));
    Odrv4 I__2302 (
            .O(N__21386),
            .I(\pwm_generator_inst.threshold_0 ));
    InMux I__2301 (
            .O(N__21383),
            .I(N__21380));
    LocalMux I__2300 (
            .O(N__21380),
            .I(N__21376));
    InMux I__2299 (
            .O(N__21379),
            .I(N__21372));
    Span4Mux_h I__2298 (
            .O(N__21376),
            .I(N__21369));
    InMux I__2297 (
            .O(N__21375),
            .I(N__21366));
    LocalMux I__2296 (
            .O(N__21372),
            .I(N__21363));
    Span4Mux_v I__2295 (
            .O(N__21369),
            .I(N__21360));
    LocalMux I__2294 (
            .O(N__21366),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__2293 (
            .O(N__21363),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__2292 (
            .O(N__21360),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2291 (
            .O(N__21353),
            .I(N__21350));
    LocalMux I__2290 (
            .O(N__21350),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__2289 (
            .O(N__21347),
            .I(N__21344));
    InMux I__2288 (
            .O(N__21344),
            .I(N__21341));
    LocalMux I__2287 (
            .O(N__21341),
            .I(N__21338));
    Odrv4 I__2286 (
            .O(N__21338),
            .I(\pwm_generator_inst.un14_counter_1 ));
    InMux I__2285 (
            .O(N__21335),
            .I(N__21332));
    LocalMux I__2284 (
            .O(N__21332),
            .I(N__21328));
    InMux I__2283 (
            .O(N__21331),
            .I(N__21324));
    Span4Mux_h I__2282 (
            .O(N__21328),
            .I(N__21321));
    InMux I__2281 (
            .O(N__21327),
            .I(N__21318));
    LocalMux I__2280 (
            .O(N__21324),
            .I(N__21315));
    Span4Mux_v I__2279 (
            .O(N__21321),
            .I(N__21312));
    LocalMux I__2278 (
            .O(N__21318),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__2277 (
            .O(N__21315),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__2276 (
            .O(N__21312),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__2275 (
            .O(N__21305),
            .I(N__21302));
    LocalMux I__2274 (
            .O(N__21302),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__2273 (
            .O(N__21299),
            .I(N__21296));
    InMux I__2272 (
            .O(N__21296),
            .I(N__21293));
    LocalMux I__2271 (
            .O(N__21293),
            .I(\pwm_generator_inst.threshold_2 ));
    InMux I__2270 (
            .O(N__21290),
            .I(N__21287));
    LocalMux I__2269 (
            .O(N__21287),
            .I(N__21284));
    Span4Mux_v I__2268 (
            .O(N__21284),
            .I(N__21279));
    InMux I__2267 (
            .O(N__21283),
            .I(N__21276));
    InMux I__2266 (
            .O(N__21282),
            .I(N__21273));
    Span4Mux_v I__2265 (
            .O(N__21279),
            .I(N__21268));
    LocalMux I__2264 (
            .O(N__21276),
            .I(N__21268));
    LocalMux I__2263 (
            .O(N__21273),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__2262 (
            .O(N__21268),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2261 (
            .O(N__21263),
            .I(N__21260));
    LocalMux I__2260 (
            .O(N__21260),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__2259 (
            .O(N__21257),
            .I(N__21254));
    LocalMux I__2258 (
            .O(N__21254),
            .I(N__21251));
    Odrv4 I__2257 (
            .O(N__21251),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    InMux I__2256 (
            .O(N__21248),
            .I(N__21245));
    LocalMux I__2255 (
            .O(N__21245),
            .I(N__21242));
    Odrv12 I__2254 (
            .O(N__21242),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8 ));
    CascadeMux I__2253 (
            .O(N__21239),
            .I(N__21235));
    CascadeMux I__2252 (
            .O(N__21238),
            .I(N__21231));
    InMux I__2251 (
            .O(N__21235),
            .I(N__21227));
    InMux I__2250 (
            .O(N__21234),
            .I(N__21224));
    InMux I__2249 (
            .O(N__21231),
            .I(N__21221));
    CascadeMux I__2248 (
            .O(N__21230),
            .I(N__21215));
    LocalMux I__2247 (
            .O(N__21227),
            .I(N__21211));
    LocalMux I__2246 (
            .O(N__21224),
            .I(N__21208));
    LocalMux I__2245 (
            .O(N__21221),
            .I(N__21205));
    CascadeMux I__2244 (
            .O(N__21220),
            .I(N__21200));
    CascadeMux I__2243 (
            .O(N__21219),
            .I(N__21197));
    InMux I__2242 (
            .O(N__21218),
            .I(N__21192));
    InMux I__2241 (
            .O(N__21215),
            .I(N__21189));
    InMux I__2240 (
            .O(N__21214),
            .I(N__21186));
    Span4Mux_v I__2239 (
            .O(N__21211),
            .I(N__21183));
    Span4Mux_v I__2238 (
            .O(N__21208),
            .I(N__21178));
    Span4Mux_v I__2237 (
            .O(N__21205),
            .I(N__21178));
    InMux I__2236 (
            .O(N__21204),
            .I(N__21165));
    InMux I__2235 (
            .O(N__21203),
            .I(N__21165));
    InMux I__2234 (
            .O(N__21200),
            .I(N__21165));
    InMux I__2233 (
            .O(N__21197),
            .I(N__21165));
    InMux I__2232 (
            .O(N__21196),
            .I(N__21165));
    InMux I__2231 (
            .O(N__21195),
            .I(N__21165));
    LocalMux I__2230 (
            .O(N__21192),
            .I(N__21158));
    LocalMux I__2229 (
            .O(N__21189),
            .I(N__21158));
    LocalMux I__2228 (
            .O(N__21186),
            .I(N__21158));
    Odrv4 I__2227 (
            .O(N__21183),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ));
    Odrv4 I__2226 (
            .O(N__21178),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ));
    LocalMux I__2225 (
            .O(N__21165),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ));
    Odrv12 I__2224 (
            .O(N__21158),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ));
    InMux I__2223 (
            .O(N__21149),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    CascadeMux I__2222 (
            .O(N__21146),
            .I(N__21143));
    InMux I__2221 (
            .O(N__21143),
            .I(N__21140));
    LocalMux I__2220 (
            .O(N__21140),
            .I(N__21136));
    InMux I__2219 (
            .O(N__21139),
            .I(N__21133));
    Sp12to4 I__2218 (
            .O(N__21136),
            .I(N__21128));
    LocalMux I__2217 (
            .O(N__21133),
            .I(N__21128));
    Odrv12 I__2216 (
            .O(N__21128),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__2215 (
            .O(N__21125),
            .I(N__21121));
    InMux I__2214 (
            .O(N__21124),
            .I(N__21117));
    LocalMux I__2213 (
            .O(N__21121),
            .I(N__21114));
    InMux I__2212 (
            .O(N__21120),
            .I(N__21111));
    LocalMux I__2211 (
            .O(N__21117),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv4 I__2210 (
            .O(N__21114),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__2209 (
            .O(N__21111),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__2208 (
            .O(N__21104),
            .I(N__21101));
    LocalMux I__2207 (
            .O(N__21101),
            .I(N__21097));
    InMux I__2206 (
            .O(N__21100),
            .I(N__21094));
    Sp12to4 I__2205 (
            .O(N__21097),
            .I(N__21089));
    LocalMux I__2204 (
            .O(N__21094),
            .I(N__21089));
    Odrv12 I__2203 (
            .O(N__21089),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8 ));
    CascadeMux I__2202 (
            .O(N__21086),
            .I(N__21083));
    InMux I__2201 (
            .O(N__21083),
            .I(N__21078));
    InMux I__2200 (
            .O(N__21082),
            .I(N__21075));
    InMux I__2199 (
            .O(N__21081),
            .I(N__21072));
    LocalMux I__2198 (
            .O(N__21078),
            .I(N__21069));
    LocalMux I__2197 (
            .O(N__21075),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__2196 (
            .O(N__21072),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    Odrv4 I__2195 (
            .O(N__21069),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    InMux I__2194 (
            .O(N__21062),
            .I(N__21058));
    InMux I__2193 (
            .O(N__21061),
            .I(N__21055));
    LocalMux I__2192 (
            .O(N__21058),
            .I(N__21052));
    LocalMux I__2191 (
            .O(N__21055),
            .I(N__21049));
    Odrv4 I__2190 (
            .O(N__21052),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8 ));
    Odrv12 I__2189 (
            .O(N__21049),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8 ));
    InMux I__2188 (
            .O(N__21044),
            .I(N__21041));
    LocalMux I__2187 (
            .O(N__21041),
            .I(N__21037));
    InMux I__2186 (
            .O(N__21040),
            .I(N__21033));
    Span4Mux_s2_h I__2185 (
            .O(N__21037),
            .I(N__21030));
    InMux I__2184 (
            .O(N__21036),
            .I(N__21027));
    LocalMux I__2183 (
            .O(N__21033),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    Odrv4 I__2182 (
            .O(N__21030),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    LocalMux I__2181 (
            .O(N__21027),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__2180 (
            .O(N__21020),
            .I(N__21017));
    LocalMux I__2179 (
            .O(N__21017),
            .I(N__21014));
    Odrv4 I__2178 (
            .O(N__21014),
            .I(un7_start_stop_0_a2));
    CascadeMux I__2177 (
            .O(N__21011),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    CascadeMux I__2176 (
            .O(N__21008),
            .I(\pwm_generator_inst.un1_counterlto9_2_cascade_ ));
    InMux I__2175 (
            .O(N__21005),
            .I(N__21002));
    LocalMux I__2174 (
            .O(N__21002),
            .I(\pwm_generator_inst.un1_counterlt9 ));
    CascadeMux I__2173 (
            .O(N__20999),
            .I(N__20996));
    InMux I__2172 (
            .O(N__20996),
            .I(N__20993));
    LocalMux I__2171 (
            .O(N__20993),
            .I(N__20990));
    Odrv4 I__2170 (
            .O(N__20990),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__2169 (
            .O(N__20987),
            .I(N__20984));
    LocalMux I__2168 (
            .O(N__20984),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791 ));
    InMux I__2167 (
            .O(N__20981),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    InMux I__2166 (
            .O(N__20978),
            .I(N__20975));
    LocalMux I__2165 (
            .O(N__20975),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    InMux I__2164 (
            .O(N__20972),
            .I(N__20969));
    LocalMux I__2163 (
            .O(N__20969),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1 ));
    InMux I__2162 (
            .O(N__20966),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__2161 (
            .O(N__20963),
            .I(N__20960));
    LocalMux I__2160 (
            .O(N__20960),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__2159 (
            .O(N__20957),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__2158 (
            .O(N__20954),
            .I(N__20951));
    LocalMux I__2157 (
            .O(N__20951),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    InMux I__2156 (
            .O(N__20948),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    InMux I__2155 (
            .O(N__20945),
            .I(N__20942));
    LocalMux I__2154 (
            .O(N__20942),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    InMux I__2153 (
            .O(N__20939),
            .I(N__20936));
    LocalMux I__2152 (
            .O(N__20936),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1 ));
    InMux I__2151 (
            .O(N__20933),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__2150 (
            .O(N__20930),
            .I(N__20927));
    LocalMux I__2149 (
            .O(N__20927),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__2148 (
            .O(N__20924),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__2147 (
            .O(N__20921),
            .I(N__20918));
    LocalMux I__2146 (
            .O(N__20918),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    InMux I__2145 (
            .O(N__20915),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    InMux I__2144 (
            .O(N__20912),
            .I(N__20909));
    LocalMux I__2143 (
            .O(N__20909),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__2142 (
            .O(N__20906),
            .I(bfn_2_18_0_));
    InMux I__2141 (
            .O(N__20903),
            .I(N__20900));
    LocalMux I__2140 (
            .O(N__20900),
            .I(N__20897));
    Odrv4 I__2139 (
            .O(N__20897),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0 ));
    InMux I__2138 (
            .O(N__20894),
            .I(N__20891));
    LocalMux I__2137 (
            .O(N__20891),
            .I(N__20888));
    Odrv4 I__2136 (
            .O(N__20888),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0 ));
    InMux I__2135 (
            .O(N__20885),
            .I(N__20882));
    LocalMux I__2134 (
            .O(N__20882),
            .I(N__20879));
    Odrv4 I__2133 (
            .O(N__20879),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0 ));
    InMux I__2132 (
            .O(N__20876),
            .I(N__20873));
    LocalMux I__2131 (
            .O(N__20873),
            .I(N__20870));
    Odrv4 I__2130 (
            .O(N__20870),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0 ));
    InMux I__2129 (
            .O(N__20867),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__2128 (
            .O(N__20864),
            .I(N__20861));
    LocalMux I__2127 (
            .O(N__20861),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__2126 (
            .O(N__20858),
            .I(N__20855));
    LocalMux I__2125 (
            .O(N__20855),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    CascadeMux I__2124 (
            .O(N__20852),
            .I(N__20849));
    InMux I__2123 (
            .O(N__20849),
            .I(N__20846));
    LocalMux I__2122 (
            .O(N__20846),
            .I(N__20843));
    Odrv4 I__2121 (
            .O(N__20843),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ));
    InMux I__2120 (
            .O(N__20840),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__2119 (
            .O(N__20837),
            .I(N__20834));
    LocalMux I__2118 (
            .O(N__20834),
            .I(N__20831));
    Odrv4 I__2117 (
            .O(N__20831),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ));
    InMux I__2116 (
            .O(N__20828),
            .I(bfn_2_15_0_));
    InMux I__2115 (
            .O(N__20825),
            .I(N__20822));
    LocalMux I__2114 (
            .O(N__20822),
            .I(N__20819));
    Odrv4 I__2113 (
            .O(N__20819),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ));
    InMux I__2112 (
            .O(N__20816),
            .I(N__20813));
    LocalMux I__2111 (
            .O(N__20813),
            .I(N__20810));
    Odrv4 I__2110 (
            .O(N__20810),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ));
    InMux I__2109 (
            .O(N__20807),
            .I(N__20804));
    LocalMux I__2108 (
            .O(N__20804),
            .I(N__20801));
    Odrv4 I__2107 (
            .O(N__20801),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ));
    InMux I__2106 (
            .O(N__20798),
            .I(N__20795));
    LocalMux I__2105 (
            .O(N__20795),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ));
    InMux I__2104 (
            .O(N__20792),
            .I(N__20789));
    LocalMux I__2103 (
            .O(N__20789),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ));
    InMux I__2102 (
            .O(N__20786),
            .I(N__20783));
    LocalMux I__2101 (
            .O(N__20783),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ));
    InMux I__2100 (
            .O(N__20780),
            .I(N__20777));
    LocalMux I__2099 (
            .O(N__20777),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ));
    CascadeMux I__2098 (
            .O(N__20774),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__2097 (
            .O(N__20771),
            .I(N__20766));
    InMux I__2096 (
            .O(N__20770),
            .I(N__20761));
    InMux I__2095 (
            .O(N__20769),
            .I(N__20761));
    LocalMux I__2094 (
            .O(N__20766),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__2093 (
            .O(N__20761),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__2092 (
            .O(N__20756),
            .I(N__20753));
    LocalMux I__2091 (
            .O(N__20753),
            .I(N__20749));
    InMux I__2090 (
            .O(N__20752),
            .I(N__20746));
    Span4Mux_v I__2089 (
            .O(N__20749),
            .I(N__20743));
    LocalMux I__2088 (
            .O(N__20746),
            .I(N__20740));
    Span4Mux_v I__2087 (
            .O(N__20743),
            .I(N__20737));
    Span4Mux_h I__2086 (
            .O(N__20740),
            .I(N__20734));
    Odrv4 I__2085 (
            .O(N__20737),
            .I(\pwm_generator_inst.un3_threshold ));
    Odrv4 I__2084 (
            .O(N__20734),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__2083 (
            .O(N__20729),
            .I(N__20726));
    LocalMux I__2082 (
            .O(N__20726),
            .I(N__20723));
    Span4Mux_h I__2081 (
            .O(N__20723),
            .I(N__20720));
    Odrv4 I__2080 (
            .O(N__20720),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__2079 (
            .O(N__20717),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__2078 (
            .O(N__20714),
            .I(N__20711));
    LocalMux I__2077 (
            .O(N__20711),
            .I(N__20708));
    Span4Mux_h I__2076 (
            .O(N__20708),
            .I(N__20705));
    Odrv4 I__2075 (
            .O(N__20705),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__2074 (
            .O(N__20702),
            .I(N__20699));
    LocalMux I__2073 (
            .O(N__20699),
            .I(N__20696));
    Span4Mux_v I__2072 (
            .O(N__20696),
            .I(N__20692));
    InMux I__2071 (
            .O(N__20695),
            .I(N__20689));
    Odrv4 I__2070 (
            .O(N__20692),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    LocalMux I__2069 (
            .O(N__20689),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    InMux I__2068 (
            .O(N__20684),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__2067 (
            .O(N__20681),
            .I(N__20678));
    LocalMux I__2066 (
            .O(N__20678),
            .I(N__20675));
    Span4Mux_h I__2065 (
            .O(N__20675),
            .I(N__20672));
    Odrv4 I__2064 (
            .O(N__20672),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__2063 (
            .O(N__20669),
            .I(N__20666));
    LocalMux I__2062 (
            .O(N__20666),
            .I(N__20662));
    InMux I__2061 (
            .O(N__20665),
            .I(N__20659));
    Odrv4 I__2060 (
            .O(N__20662),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    LocalMux I__2059 (
            .O(N__20659),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    InMux I__2058 (
            .O(N__20654),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__2057 (
            .O(N__20651),
            .I(N__20648));
    LocalMux I__2056 (
            .O(N__20648),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__2055 (
            .O(N__20645),
            .I(N__20642));
    LocalMux I__2054 (
            .O(N__20642),
            .I(N__20638));
    InMux I__2053 (
            .O(N__20641),
            .I(N__20635));
    Odrv4 I__2052 (
            .O(N__20638),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    LocalMux I__2051 (
            .O(N__20635),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    InMux I__2050 (
            .O(N__20630),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    CascadeMux I__2049 (
            .O(N__20627),
            .I(N__20624));
    InMux I__2048 (
            .O(N__20624),
            .I(N__20621));
    LocalMux I__2047 (
            .O(N__20621),
            .I(N__20618));
    Odrv4 I__2046 (
            .O(N__20618),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ));
    InMux I__2045 (
            .O(N__20615),
            .I(N__20612));
    LocalMux I__2044 (
            .O(N__20612),
            .I(N__20608));
    InMux I__2043 (
            .O(N__20611),
            .I(N__20605));
    Odrv4 I__2042 (
            .O(N__20608),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8 ));
    LocalMux I__2041 (
            .O(N__20605),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8 ));
    InMux I__2040 (
            .O(N__20600),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__2039 (
            .O(N__20597),
            .I(N__20594));
    LocalMux I__2038 (
            .O(N__20594),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ));
    InMux I__2037 (
            .O(N__20591),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__2036 (
            .O(N__20588),
            .I(N__20585));
    LocalMux I__2035 (
            .O(N__20585),
            .I(N__20580));
    InMux I__2034 (
            .O(N__20584),
            .I(N__20575));
    InMux I__2033 (
            .O(N__20583),
            .I(N__20575));
    Span4Mux_s2_h I__2032 (
            .O(N__20580),
            .I(N__20572));
    LocalMux I__2031 (
            .O(N__20575),
            .I(pwm_duty_input_6));
    Odrv4 I__2030 (
            .O(N__20572),
            .I(pwm_duty_input_6));
    InMux I__2029 (
            .O(N__20567),
            .I(N__20560));
    InMux I__2028 (
            .O(N__20566),
            .I(N__20560));
    InMux I__2027 (
            .O(N__20565),
            .I(N__20557));
    LocalMux I__2026 (
            .O(N__20560),
            .I(pwm_duty_input_8));
    LocalMux I__2025 (
            .O(N__20557),
            .I(pwm_duty_input_8));
    CascadeMux I__2024 (
            .O(N__20552),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__2023 (
            .O(N__20549),
            .I(N__20545));
    CascadeMux I__2022 (
            .O(N__20548),
            .I(N__20541));
    LocalMux I__2021 (
            .O(N__20545),
            .I(N__20538));
    InMux I__2020 (
            .O(N__20544),
            .I(N__20533));
    InMux I__2019 (
            .O(N__20541),
            .I(N__20533));
    Span4Mux_s1_h I__2018 (
            .O(N__20538),
            .I(N__20530));
    LocalMux I__2017 (
            .O(N__20533),
            .I(pwm_duty_input_9));
    Odrv4 I__2016 (
            .O(N__20530),
            .I(pwm_duty_input_9));
    InMux I__2015 (
            .O(N__20525),
            .I(N__20522));
    LocalMux I__2014 (
            .O(N__20522),
            .I(N__20517));
    InMux I__2013 (
            .O(N__20521),
            .I(N__20514));
    InMux I__2012 (
            .O(N__20520),
            .I(N__20511));
    Span4Mux_s1_h I__2011 (
            .O(N__20517),
            .I(N__20508));
    LocalMux I__2010 (
            .O(N__20514),
            .I(pwm_duty_input_3));
    LocalMux I__2009 (
            .O(N__20511),
            .I(pwm_duty_input_3));
    Odrv4 I__2008 (
            .O(N__20508),
            .I(pwm_duty_input_3));
    CascadeMux I__2007 (
            .O(N__20501),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ));
    InMux I__2006 (
            .O(N__20498),
            .I(N__20495));
    LocalMux I__2005 (
            .O(N__20495),
            .I(N__20490));
    InMux I__2004 (
            .O(N__20494),
            .I(N__20487));
    InMux I__2003 (
            .O(N__20493),
            .I(N__20484));
    Span4Mux_v I__2002 (
            .O(N__20490),
            .I(N__20481));
    LocalMux I__2001 (
            .O(N__20487),
            .I(pwm_duty_input_4));
    LocalMux I__2000 (
            .O(N__20484),
            .I(pwm_duty_input_4));
    Odrv4 I__1999 (
            .O(N__20481),
            .I(pwm_duty_input_4));
    InMux I__1998 (
            .O(N__20474),
            .I(N__20471));
    LocalMux I__1997 (
            .O(N__20471),
            .I(N__20467));
    InMux I__1996 (
            .O(N__20470),
            .I(N__20464));
    Span4Mux_s1_h I__1995 (
            .O(N__20467),
            .I(N__20461));
    LocalMux I__1994 (
            .O(N__20464),
            .I(pwm_duty_input_0));
    Odrv4 I__1993 (
            .O(N__20461),
            .I(pwm_duty_input_0));
    InMux I__1992 (
            .O(N__20456),
            .I(N__20452));
    InMux I__1991 (
            .O(N__20455),
            .I(N__20449));
    LocalMux I__1990 (
            .O(N__20452),
            .I(pwm_duty_input_1));
    LocalMux I__1989 (
            .O(N__20449),
            .I(pwm_duty_input_1));
    InMux I__1988 (
            .O(N__20444),
            .I(N__20440));
    InMux I__1987 (
            .O(N__20443),
            .I(N__20437));
    LocalMux I__1986 (
            .O(N__20440),
            .I(pwm_duty_input_2));
    LocalMux I__1985 (
            .O(N__20437),
            .I(pwm_duty_input_2));
    InMux I__1984 (
            .O(N__20432),
            .I(N__20429));
    LocalMux I__1983 (
            .O(N__20429),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__1982 (
            .O(N__20426),
            .I(N__20423));
    LocalMux I__1981 (
            .O(N__20423),
            .I(N__20420));
    Odrv4 I__1980 (
            .O(N__20420),
            .I(\current_shift_inst.PI_CTRL.N_140 ));
    InMux I__1979 (
            .O(N__20417),
            .I(N__20414));
    LocalMux I__1978 (
            .O(N__20414),
            .I(N__20411));
    Odrv4 I__1977 (
            .O(N__20411),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    CascadeMux I__1976 (
            .O(N__20408),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_ ));
    CascadeMux I__1975 (
            .O(N__20405),
            .I(N__20400));
    CascadeMux I__1974 (
            .O(N__20404),
            .I(N__20397));
    CascadeMux I__1973 (
            .O(N__20403),
            .I(N__20394));
    InMux I__1972 (
            .O(N__20400),
            .I(N__20391));
    InMux I__1971 (
            .O(N__20397),
            .I(N__20386));
    InMux I__1970 (
            .O(N__20394),
            .I(N__20386));
    LocalMux I__1969 (
            .O(N__20391),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    LocalMux I__1968 (
            .O(N__20386),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1967 (
            .O(N__20381),
            .I(N__20372));
    InMux I__1966 (
            .O(N__20380),
            .I(N__20372));
    InMux I__1965 (
            .O(N__20379),
            .I(N__20372));
    LocalMux I__1964 (
            .O(N__20372),
            .I(N__20369));
    Odrv4 I__1963 (
            .O(N__20369),
            .I(\current_shift_inst.PI_CTRL.N_145 ));
    InMux I__1962 (
            .O(N__20366),
            .I(N__20363));
    LocalMux I__1961 (
            .O(N__20363),
            .I(N__20358));
    InMux I__1960 (
            .O(N__20362),
            .I(N__20355));
    InMux I__1959 (
            .O(N__20361),
            .I(N__20352));
    Span4Mux_v I__1958 (
            .O(N__20358),
            .I(N__20349));
    LocalMux I__1957 (
            .O(N__20355),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__1956 (
            .O(N__20352),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    Odrv4 I__1955 (
            .O(N__20349),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    CascadeMux I__1954 (
            .O(N__20342),
            .I(N__20339));
    InMux I__1953 (
            .O(N__20339),
            .I(N__20336));
    LocalMux I__1952 (
            .O(N__20336),
            .I(N__20333));
    Odrv12 I__1951 (
            .O(N__20333),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__1950 (
            .O(N__20330),
            .I(bfn_1_21_0_));
    InMux I__1949 (
            .O(N__20327),
            .I(N__20324));
    LocalMux I__1948 (
            .O(N__20324),
            .I(N__20321));
    Odrv12 I__1947 (
            .O(N__20321),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__1946 (
            .O(N__20318),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__1945 (
            .O(N__20315),
            .I(N__20312));
    LocalMux I__1944 (
            .O(N__20312),
            .I(N__20309));
    Odrv4 I__1943 (
            .O(N__20309),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__1942 (
            .O(N__20306),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__1941 (
            .O(N__20303),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__1940 (
            .O(N__20300),
            .I(N__20297));
    LocalMux I__1939 (
            .O(N__20297),
            .I(N_42_i_i));
    InMux I__1938 (
            .O(N__20294),
            .I(N__20291));
    LocalMux I__1937 (
            .O(N__20291),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    InMux I__1936 (
            .O(N__20288),
            .I(N__20281));
    InMux I__1935 (
            .O(N__20287),
            .I(N__20281));
    InMux I__1934 (
            .O(N__20286),
            .I(N__20278));
    LocalMux I__1933 (
            .O(N__20281),
            .I(pwm_duty_input_7));
    LocalMux I__1932 (
            .O(N__20278),
            .I(pwm_duty_input_7));
    InMux I__1931 (
            .O(N__20273),
            .I(N__20269));
    CascadeMux I__1930 (
            .O(N__20272),
            .I(N__20266));
    LocalMux I__1929 (
            .O(N__20269),
            .I(N__20262));
    InMux I__1928 (
            .O(N__20266),
            .I(N__20259));
    InMux I__1927 (
            .O(N__20265),
            .I(N__20256));
    Span4Mux_s1_h I__1926 (
            .O(N__20262),
            .I(N__20253));
    LocalMux I__1925 (
            .O(N__20259),
            .I(pwm_duty_input_5));
    LocalMux I__1924 (
            .O(N__20256),
            .I(pwm_duty_input_5));
    Odrv4 I__1923 (
            .O(N__20253),
            .I(pwm_duty_input_5));
    InMux I__1922 (
            .O(N__20246),
            .I(N__20243));
    LocalMux I__1921 (
            .O(N__20243),
            .I(N__20240));
    Span4Mux_v I__1920 (
            .O(N__20240),
            .I(N__20237));
    Span4Mux_v I__1919 (
            .O(N__20237),
            .I(N__20234));
    Odrv4 I__1918 (
            .O(N__20234),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1917 (
            .O(N__20231),
            .I(N__20228));
    LocalMux I__1916 (
            .O(N__20228),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__1915 (
            .O(N__20225),
            .I(N__20222));
    LocalMux I__1914 (
            .O(N__20222),
            .I(N__20219));
    Span12Mux_h I__1913 (
            .O(N__20219),
            .I(N__20216));
    Odrv12 I__1912 (
            .O(N__20216),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1911 (
            .O(N__20213),
            .I(N__20210));
    LocalMux I__1910 (
            .O(N__20210),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__1909 (
            .O(N__20207),
            .I(N__20204));
    LocalMux I__1908 (
            .O(N__20204),
            .I(N__20200));
    InMux I__1907 (
            .O(N__20203),
            .I(N__20197));
    Span4Mux_v I__1906 (
            .O(N__20200),
            .I(N__20194));
    LocalMux I__1905 (
            .O(N__20197),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__1904 (
            .O(N__20194),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    InMux I__1903 (
            .O(N__20189),
            .I(N__20186));
    LocalMux I__1902 (
            .O(N__20186),
            .I(N__20183));
    Odrv12 I__1901 (
            .O(N__20183),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    InMux I__1900 (
            .O(N__20180),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    InMux I__1899 (
            .O(N__20177),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    InMux I__1898 (
            .O(N__20174),
            .I(N__20171));
    LocalMux I__1897 (
            .O(N__20171),
            .I(N__20168));
    Odrv12 I__1896 (
            .O(N__20168),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    InMux I__1895 (
            .O(N__20165),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__1894 (
            .O(N__20162),
            .I(N__20157));
    InMux I__1893 (
            .O(N__20161),
            .I(N__20154));
    InMux I__1892 (
            .O(N__20160),
            .I(N__20151));
    LocalMux I__1891 (
            .O(N__20157),
            .I(N__20148));
    LocalMux I__1890 (
            .O(N__20154),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    LocalMux I__1889 (
            .O(N__20151),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    Odrv12 I__1888 (
            .O(N__20148),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    InMux I__1887 (
            .O(N__20141),
            .I(N__20138));
    LocalMux I__1886 (
            .O(N__20138),
            .I(N__20135));
    Odrv12 I__1885 (
            .O(N__20135),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    InMux I__1884 (
            .O(N__20132),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__1883 (
            .O(N__20129),
            .I(N__20124));
    InMux I__1882 (
            .O(N__20128),
            .I(N__20121));
    InMux I__1881 (
            .O(N__20127),
            .I(N__20118));
    LocalMux I__1880 (
            .O(N__20124),
            .I(N__20115));
    LocalMux I__1879 (
            .O(N__20121),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    LocalMux I__1878 (
            .O(N__20118),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv12 I__1877 (
            .O(N__20115),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__1876 (
            .O(N__20108),
            .I(N__20105));
    LocalMux I__1875 (
            .O(N__20105),
            .I(N__20102));
    Span4Mux_h I__1874 (
            .O(N__20102),
            .I(N__20099));
    Span4Mux_v I__1873 (
            .O(N__20099),
            .I(N__20096));
    Odrv4 I__1872 (
            .O(N__20096),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    InMux I__1871 (
            .O(N__20093),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    CascadeMux I__1870 (
            .O(N__20090),
            .I(N__20086));
    CascadeMux I__1869 (
            .O(N__20089),
            .I(N__20082));
    InMux I__1868 (
            .O(N__20086),
            .I(N__20079));
    InMux I__1867 (
            .O(N__20085),
            .I(N__20076));
    InMux I__1866 (
            .O(N__20082),
            .I(N__20073));
    LocalMux I__1865 (
            .O(N__20079),
            .I(N__20070));
    LocalMux I__1864 (
            .O(N__20076),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__1863 (
            .O(N__20073),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    Odrv12 I__1862 (
            .O(N__20070),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    InMux I__1861 (
            .O(N__20063),
            .I(N__20060));
    LocalMux I__1860 (
            .O(N__20060),
            .I(N__20057));
    Odrv12 I__1859 (
            .O(N__20057),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    InMux I__1858 (
            .O(N__20054),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    InMux I__1857 (
            .O(N__20051),
            .I(N__20048));
    LocalMux I__1856 (
            .O(N__20048),
            .I(N__20045));
    Span4Mux_v I__1855 (
            .O(N__20045),
            .I(N__20042));
    Span4Mux_v I__1854 (
            .O(N__20042),
            .I(N__20039));
    Odrv4 I__1853 (
            .O(N__20039),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1852 (
            .O(N__20036),
            .I(N__20033));
    LocalMux I__1851 (
            .O(N__20033),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__1850 (
            .O(N__20030),
            .I(N__20027));
    LocalMux I__1849 (
            .O(N__20027),
            .I(N__20024));
    Span12Mux_h I__1848 (
            .O(N__20024),
            .I(N__20021));
    Odrv12 I__1847 (
            .O(N__20021),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1846 (
            .O(N__20018),
            .I(N__20015));
    LocalMux I__1845 (
            .O(N__20015),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__1844 (
            .O(N__20012),
            .I(N__20009));
    LocalMux I__1843 (
            .O(N__20009),
            .I(N__20006));
    Span4Mux_v I__1842 (
            .O(N__20006),
            .I(N__20003));
    Span4Mux_v I__1841 (
            .O(N__20003),
            .I(N__20000));
    Odrv4 I__1840 (
            .O(N__20000),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1839 (
            .O(N__19997),
            .I(N__19994));
    LocalMux I__1838 (
            .O(N__19994),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__1837 (
            .O(N__19991),
            .I(N__19988));
    LocalMux I__1836 (
            .O(N__19988),
            .I(N__19985));
    Span4Mux_v I__1835 (
            .O(N__19985),
            .I(N__19982));
    Span4Mux_v I__1834 (
            .O(N__19982),
            .I(N__19979));
    Span4Mux_v I__1833 (
            .O(N__19979),
            .I(N__19976));
    Odrv4 I__1832 (
            .O(N__19976),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1831 (
            .O(N__19973),
            .I(N__19970));
    LocalMux I__1830 (
            .O(N__19970),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__1829 (
            .O(N__19967),
            .I(N__19964));
    LocalMux I__1828 (
            .O(N__19964),
            .I(N__19961));
    Span4Mux_v I__1827 (
            .O(N__19961),
            .I(N__19958));
    Span4Mux_v I__1826 (
            .O(N__19958),
            .I(N__19955));
    Odrv4 I__1825 (
            .O(N__19955),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1824 (
            .O(N__19952),
            .I(N__19949));
    LocalMux I__1823 (
            .O(N__19949),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    InMux I__1822 (
            .O(N__19946),
            .I(N__19943));
    LocalMux I__1821 (
            .O(N__19943),
            .I(N__19940));
    Span4Mux_v I__1820 (
            .O(N__19940),
            .I(N__19937));
    Span4Mux_v I__1819 (
            .O(N__19937),
            .I(N__19934));
    Odrv4 I__1818 (
            .O(N__19934),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1817 (
            .O(N__19931),
            .I(N__19928));
    LocalMux I__1816 (
            .O(N__19928),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__1815 (
            .O(N__19925),
            .I(N__19922));
    LocalMux I__1814 (
            .O(N__19922),
            .I(N__19919));
    Span4Mux_v I__1813 (
            .O(N__19919),
            .I(N__19916));
    Span4Mux_v I__1812 (
            .O(N__19916),
            .I(N__19913));
    Odrv4 I__1811 (
            .O(N__19913),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1810 (
            .O(N__19910),
            .I(N__19907));
    LocalMux I__1809 (
            .O(N__19907),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__1808 (
            .O(N__19904),
            .I(N__19901));
    LocalMux I__1807 (
            .O(N__19901),
            .I(N__19898));
    Span4Mux_v I__1806 (
            .O(N__19898),
            .I(N__19895));
    Span4Mux_v I__1805 (
            .O(N__19895),
            .I(N__19892));
    Odrv4 I__1804 (
            .O(N__19892),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1803 (
            .O(N__19889),
            .I(N__19886));
    LocalMux I__1802 (
            .O(N__19886),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__1801 (
            .O(N__19883),
            .I(N__19877));
    InMux I__1800 (
            .O(N__19882),
            .I(N__19877));
    LocalMux I__1799 (
            .O(N__19877),
            .I(N__19874));
    Span4Mux_v I__1798 (
            .O(N__19874),
            .I(N__19871));
    Odrv4 I__1797 (
            .O(N__19871),
            .I(\pwm_generator_inst.O_10 ));
    CascadeMux I__1796 (
            .O(N__19868),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10_cascade_ ));
    CascadeMux I__1795 (
            .O(N__19865),
            .I(N__19862));
    InMux I__1794 (
            .O(N__19862),
            .I(N__19859));
    LocalMux I__1793 (
            .O(N__19859),
            .I(N__19856));
    Span4Mux_v I__1792 (
            .O(N__19856),
            .I(N__19853));
    Span4Mux_v I__1791 (
            .O(N__19853),
            .I(N__19850));
    Odrv4 I__1790 (
            .O(N__19850),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__1789 (
            .O(N__19847),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    CascadeMux I__1788 (
            .O(N__19844),
            .I(N__19841));
    InMux I__1787 (
            .O(N__19841),
            .I(N__19838));
    LocalMux I__1786 (
            .O(N__19838),
            .I(N__19835));
    Span4Mux_v I__1785 (
            .O(N__19835),
            .I(N__19832));
    Span4Mux_v I__1784 (
            .O(N__19832),
            .I(N__19829));
    Odrv4 I__1783 (
            .O(N__19829),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    InMux I__1782 (
            .O(N__19826),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    CascadeMux I__1781 (
            .O(N__19823),
            .I(N__19820));
    InMux I__1780 (
            .O(N__19820),
            .I(N__19817));
    LocalMux I__1779 (
            .O(N__19817),
            .I(N__19814));
    Span4Mux_v I__1778 (
            .O(N__19814),
            .I(N__19811));
    Span4Mux_v I__1777 (
            .O(N__19811),
            .I(N__19808));
    Odrv4 I__1776 (
            .O(N__19808),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__1775 (
            .O(N__19805),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    InMux I__1774 (
            .O(N__19802),
            .I(N__19796));
    InMux I__1773 (
            .O(N__19801),
            .I(N__19796));
    LocalMux I__1772 (
            .O(N__19796),
            .I(N__19793));
    Span4Mux_v I__1771 (
            .O(N__19793),
            .I(N__19784));
    InMux I__1770 (
            .O(N__19792),
            .I(N__19777));
    InMux I__1769 (
            .O(N__19791),
            .I(N__19777));
    InMux I__1768 (
            .O(N__19790),
            .I(N__19777));
    InMux I__1767 (
            .O(N__19789),
            .I(N__19770));
    InMux I__1766 (
            .O(N__19788),
            .I(N__19770));
    InMux I__1765 (
            .O(N__19787),
            .I(N__19770));
    Odrv4 I__1764 (
            .O(N__19784),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    LocalMux I__1763 (
            .O(N__19777),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    LocalMux I__1762 (
            .O(N__19770),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    CascadeMux I__1761 (
            .O(N__19763),
            .I(N__19760));
    InMux I__1760 (
            .O(N__19760),
            .I(N__19757));
    LocalMux I__1759 (
            .O(N__19757),
            .I(N__19754));
    Odrv12 I__1758 (
            .O(N__19754),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    InMux I__1757 (
            .O(N__19751),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__1756 (
            .O(N__19748),
            .I(N__19745));
    LocalMux I__1755 (
            .O(N__19745),
            .I(N__19742));
    Span12Mux_v I__1754 (
            .O(N__19742),
            .I(N__19739));
    Odrv12 I__1753 (
            .O(N__19739),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__1752 (
            .O(N__19736),
            .I(bfn_1_15_0_));
    InMux I__1751 (
            .O(N__19733),
            .I(N__19730));
    LocalMux I__1750 (
            .O(N__19730),
            .I(N__19727));
    Span4Mux_v I__1749 (
            .O(N__19727),
            .I(N__19724));
    Span4Mux_v I__1748 (
            .O(N__19724),
            .I(N__19721));
    Odrv4 I__1747 (
            .O(N__19721),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    CascadeMux I__1746 (
            .O(N__19718),
            .I(N__19715));
    InMux I__1745 (
            .O(N__19715),
            .I(N__19712));
    LocalMux I__1744 (
            .O(N__19712),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__1743 (
            .O(N__19709),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__1742 (
            .O(N__19706),
            .I(N__19703));
    LocalMux I__1741 (
            .O(N__19703),
            .I(N__19700));
    Span4Mux_v I__1740 (
            .O(N__19700),
            .I(N__19697));
    Span4Mux_v I__1739 (
            .O(N__19697),
            .I(N__19694));
    Odrv4 I__1738 (
            .O(N__19694),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__1737 (
            .O(N__19691),
            .I(N__19688));
    InMux I__1736 (
            .O(N__19688),
            .I(N__19685));
    LocalMux I__1735 (
            .O(N__19685),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    InMux I__1734 (
            .O(N__19682),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__1733 (
            .O(N__19679),
            .I(N__19676));
    LocalMux I__1732 (
            .O(N__19676),
            .I(N__19673));
    Span4Mux_v I__1731 (
            .O(N__19673),
            .I(N__19670));
    Span4Mux_v I__1730 (
            .O(N__19670),
            .I(N__19667));
    Odrv4 I__1729 (
            .O(N__19667),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    CascadeMux I__1728 (
            .O(N__19664),
            .I(N__19661));
    InMux I__1727 (
            .O(N__19661),
            .I(N__19658));
    LocalMux I__1726 (
            .O(N__19658),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    InMux I__1725 (
            .O(N__19655),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__1724 (
            .O(N__19652),
            .I(N__19649));
    LocalMux I__1723 (
            .O(N__19649),
            .I(N__19646));
    Span4Mux_v I__1722 (
            .O(N__19646),
            .I(N__19643));
    Span4Mux_v I__1721 (
            .O(N__19643),
            .I(N__19640));
    Odrv4 I__1720 (
            .O(N__19640),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    CascadeMux I__1719 (
            .O(N__19637),
            .I(N__19634));
    InMux I__1718 (
            .O(N__19634),
            .I(N__19631));
    LocalMux I__1717 (
            .O(N__19631),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    InMux I__1716 (
            .O(N__19628),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__1715 (
            .O(N__19625),
            .I(N__19622));
    LocalMux I__1714 (
            .O(N__19622),
            .I(N__19619));
    Span12Mux_h I__1713 (
            .O(N__19619),
            .I(N__19616));
    Odrv12 I__1712 (
            .O(N__19616),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    CascadeMux I__1711 (
            .O(N__19613),
            .I(N__19610));
    InMux I__1710 (
            .O(N__19610),
            .I(N__19607));
    LocalMux I__1709 (
            .O(N__19607),
            .I(N__19604));
    Span4Mux_h I__1708 (
            .O(N__19604),
            .I(N__19601));
    Odrv4 I__1707 (
            .O(N__19601),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    InMux I__1706 (
            .O(N__19598),
            .I(bfn_1_14_0_));
    InMux I__1705 (
            .O(N__19595),
            .I(N__19592));
    LocalMux I__1704 (
            .O(N__19592),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    CascadeMux I__1703 (
            .O(N__19589),
            .I(N__19586));
    InMux I__1702 (
            .O(N__19586),
            .I(N__19583));
    LocalMux I__1701 (
            .O(N__19583),
            .I(N__19580));
    Span4Mux_v I__1700 (
            .O(N__19580),
            .I(N__19577));
    Span4Mux_v I__1699 (
            .O(N__19577),
            .I(N__19574));
    Odrv4 I__1698 (
            .O(N__19574),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    InMux I__1697 (
            .O(N__19571),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    CascadeMux I__1696 (
            .O(N__19568),
            .I(N__19565));
    InMux I__1695 (
            .O(N__19565),
            .I(N__19562));
    LocalMux I__1694 (
            .O(N__19562),
            .I(N__19559));
    Span4Mux_v I__1693 (
            .O(N__19559),
            .I(N__19556));
    Span4Mux_v I__1692 (
            .O(N__19556),
            .I(N__19553));
    Odrv4 I__1691 (
            .O(N__19553),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__1690 (
            .O(N__19550),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    CascadeMux I__1689 (
            .O(N__19547),
            .I(N__19544));
    InMux I__1688 (
            .O(N__19544),
            .I(N__19541));
    LocalMux I__1687 (
            .O(N__19541),
            .I(N__19538));
    Span4Mux_v I__1686 (
            .O(N__19538),
            .I(N__19535));
    Span4Mux_v I__1685 (
            .O(N__19535),
            .I(N__19532));
    Odrv4 I__1684 (
            .O(N__19532),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__1683 (
            .O(N__19529),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    InMux I__1682 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__1681 (
            .O(N__19523),
            .I(N__19520));
    Span12Mux_h I__1680 (
            .O(N__19520),
            .I(N__19517));
    Odrv12 I__1679 (
            .O(N__19517),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__1678 (
            .O(N__19514),
            .I(N__19511));
    InMux I__1677 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__1676 (
            .O(N__19508),
            .I(N__19505));
    Span4Mux_h I__1675 (
            .O(N__19505),
            .I(N__19502));
    Odrv4 I__1674 (
            .O(N__19502),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__1673 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__1672 (
            .O(N__19496),
            .I(N__19493));
    Span4Mux_v I__1671 (
            .O(N__19493),
            .I(N__19490));
    Span4Mux_v I__1670 (
            .O(N__19490),
            .I(N__19487));
    Odrv4 I__1669 (
            .O(N__19487),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__1668 (
            .O(N__19484),
            .I(N__19481));
    InMux I__1667 (
            .O(N__19481),
            .I(N__19478));
    LocalMux I__1666 (
            .O(N__19478),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    InMux I__1665 (
            .O(N__19475),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__1664 (
            .O(N__19472),
            .I(N__19469));
    LocalMux I__1663 (
            .O(N__19469),
            .I(N__19466));
    Span4Mux_v I__1662 (
            .O(N__19466),
            .I(N__19463));
    Span4Mux_v I__1661 (
            .O(N__19463),
            .I(N__19460));
    Odrv4 I__1660 (
            .O(N__19460),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__1659 (
            .O(N__19457),
            .I(N__19454));
    InMux I__1658 (
            .O(N__19454),
            .I(N__19451));
    LocalMux I__1657 (
            .O(N__19451),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__1656 (
            .O(N__19448),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__1655 (
            .O(N__19445),
            .I(N__19442));
    LocalMux I__1654 (
            .O(N__19442),
            .I(N__19439));
    Span4Mux_v I__1653 (
            .O(N__19439),
            .I(N__19436));
    Span4Mux_v I__1652 (
            .O(N__19436),
            .I(N__19433));
    Odrv4 I__1651 (
            .O(N__19433),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__1650 (
            .O(N__19430),
            .I(N__19427));
    InMux I__1649 (
            .O(N__19427),
            .I(N__19424));
    LocalMux I__1648 (
            .O(N__19424),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    InMux I__1647 (
            .O(N__19421),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__1646 (
            .O(N__19418),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__1645 (
            .O(N__19415),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__1644 (
            .O(N__19412),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__1643 (
            .O(N__19409),
            .I(bfn_1_10_0_));
    InMux I__1642 (
            .O(N__19406),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__1641 (
            .O(N__19403),
            .I(N__19400));
    LocalMux I__1640 (
            .O(N__19400),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__1639 (
            .O(N__19397),
            .I(N__19391));
    InMux I__1638 (
            .O(N__19396),
            .I(N__19391));
    LocalMux I__1637 (
            .O(N__19391),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    InMux I__1636 (
            .O(N__19388),
            .I(bfn_1_9_0_));
    InMux I__1635 (
            .O(N__19385),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__1634 (
            .O(N__19382),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__1633 (
            .O(N__19379),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__1632 (
            .O(N__19376),
            .I(\pwm_generator_inst.counter_cry_3 ));
    IoInMux I__1631 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__1630 (
            .O(N__19370),
            .I(N__19367));
    Span4Mux_s3_v I__1629 (
            .O(N__19367),
            .I(N__19364));
    Span4Mux_h I__1628 (
            .O(N__19364),
            .I(N__19361));
    Sp12to4 I__1627 (
            .O(N__19361),
            .I(N__19358));
    Span12Mux_s9_v I__1626 (
            .O(N__19358),
            .I(N__19355));
    Span12Mux_v I__1625 (
            .O(N__19355),
            .I(N__19352));
    Odrv12 I__1624 (
            .O(N__19352),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1623 (
            .O(N__19349),
            .I(N__19346));
    LocalMux I__1622 (
            .O(N__19346),
            .I(N__19343));
    IoSpan4Mux I__1621 (
            .O(N__19343),
            .I(N__19340));
    IoSpan4Mux I__1620 (
            .O(N__19340),
            .I(N__19337));
    Odrv4 I__1619 (
            .O(N__19337),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_18_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_7_0_));
    defparam IN_MUX_bfv_18_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_8_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_18_8_0_));
    defparam IN_MUX_bfv_18_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_9_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_18_9_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_1_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_21_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_1_21_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_5_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_5_16_0_));
    defparam IN_MUX_bfv_5_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_17_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_5_17_0_));
    defparam IN_MUX_bfv_5_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_5_18_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_12_14_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19373),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19349),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__35582),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_167_i_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__24037),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un1_start_g ));
    ICE_GB \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0  (
            .USERSIGNALTOGLOBALBUFFER(N__37436),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_hc.un1_start_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__45040),
            .CLKHFEN(N__45044),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__45088),
            .RGB2PWM(N__20300),
            .RGB1(rgb_g),
            .CURREN(N__45045),
            .RGB2(rgb_b),
            .RGB1PWM(N__21020),
            .RGB0PWM(N__48683),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_5_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23198),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49148),
            .ce(),
            .sr(N__48597));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_6_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_6_0 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_6_0  (
            .in0(N__19397),
            .in1(N__19403),
            .in2(N__21968),
            .in3(N__19801),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_2  (
            .in0(N__19396),
            .in1(N__21924),
            .in2(_gnd_net_),
            .in3(N__19802),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_1_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_1_9_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_1_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_1_9_0  (
            .in0(N__21518),
            .in1(N__21375),
            .in2(_gnd_net_),
            .in3(N__19388),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__49147),
            .ce(),
            .sr(N__48629));
    defparam \pwm_generator_inst.counter_1_LC_1_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_1_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_1_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_1_9_1  (
            .in0(N__21514),
            .in1(N__21327),
            .in2(_gnd_net_),
            .in3(N__19385),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__49147),
            .ce(),
            .sr(N__48629));
    defparam \pwm_generator_inst.counter_2_LC_1_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_1_9_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_1_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_1_9_2  (
            .in0(N__21519),
            .in1(N__21282),
            .in2(_gnd_net_),
            .in3(N__19382),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__49147),
            .ce(),
            .sr(N__48629));
    defparam \pwm_generator_inst.counter_3_LC_1_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_1_9_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_1_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_1_9_3  (
            .in0(N__21515),
            .in1(N__21795),
            .in2(_gnd_net_),
            .in3(N__19379),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__49147),
            .ce(),
            .sr(N__48629));
    defparam \pwm_generator_inst.counter_4_LC_1_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_1_9_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_1_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_1_9_4  (
            .in0(N__21520),
            .in1(N__21753),
            .in2(_gnd_net_),
            .in3(N__19376),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__49147),
            .ce(),
            .sr(N__48629));
    defparam \pwm_generator_inst.counter_5_LC_1_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_1_9_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_1_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_1_9_5  (
            .in0(N__21516),
            .in1(N__21702),
            .in2(_gnd_net_),
            .in3(N__19418),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__49147),
            .ce(),
            .sr(N__48629));
    defparam \pwm_generator_inst.counter_6_LC_1_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_1_9_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_1_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_1_9_6  (
            .in0(N__21521),
            .in1(N__21654),
            .in2(_gnd_net_),
            .in3(N__19415),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__49147),
            .ce(),
            .sr(N__48629));
    defparam \pwm_generator_inst.counter_7_LC_1_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_1_9_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_1_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_1_9_7  (
            .in0(N__21517),
            .in1(N__21618),
            .in2(_gnd_net_),
            .in3(N__19412),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__49147),
            .ce(),
            .sr(N__48629));
    defparam \pwm_generator_inst.counter_8_LC_1_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_1_10_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_1_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_1_10_0  (
            .in0(N__21513),
            .in1(N__21586),
            .in2(_gnd_net_),
            .in3(N__19409),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__49146),
            .ce(),
            .sr(N__48636));
    defparam \pwm_generator_inst.counter_9_LC_1_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_1_10_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_1_10_1  (
            .in0(N__21549),
            .in1(N__21512),
            .in2(_gnd_net_),
            .in3(N__19406),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49146),
            .ce(),
            .sr(N__48636));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3  (
            .in0(N__22404),
            .in1(N__22711),
            .in2(N__21824),
            .in3(N__20426),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49146),
            .ce(),
            .sr(N__48636));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_4 .LUT_INIT=16'b1000100011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_4  (
            .in0(N__22658),
            .in1(N__22405),
            .in2(N__22303),
            .in3(N__23190),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49146),
            .ce(),
            .sr(N__48636));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_6 .LUT_INIT=16'b1000100011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_6  (
            .in0(N__22961),
            .in1(N__22406),
            .in2(N__22304),
            .in3(N__23191),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49146),
            .ce(),
            .sr(N__48636));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7  (
            .in0(N__22295),
            .in1(N__20417),
            .in2(N__22760),
            .in3(N__21473),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49146),
            .ce(),
            .sr(N__48636));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0  (
            .in0(N__21471),
            .in1(N__22775),
            .in2(N__20404),
            .in3(N__20381),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49144),
            .ce(),
            .sr(N__48639));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_1 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_1  (
            .in0(N__20379),
            .in1(N__22505),
            .in2(N__20405),
            .in3(N__21472),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49144),
            .ce(),
            .sr(N__48639));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_11_5 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_11_5  (
            .in0(N__23189),
            .in1(N__22294),
            .in2(N__22571),
            .in3(N__22407),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49144),
            .ce(),
            .sr(N__48639));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_11_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_11_6  (
            .in0(N__21470),
            .in1(N__22796),
            .in2(N__20403),
            .in3(N__20380),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49144),
            .ce(),
            .sr(N__48639));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4 .LUT_INIT=16'b1010000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4  (
            .in0(N__22537),
            .in1(N__22293),
            .in2(N__22408),
            .in3(N__23187),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49141),
            .ce(),
            .sr(N__48643));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_1_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_1_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__19526),
            .in2(N__19514),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__19499),
            .in2(N__19484),
            .in3(N__19475),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__19472),
            .in2(N__19457),
            .in3(N__19448),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__19445),
            .in2(N__19430),
            .in3(N__19421),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__19733),
            .in2(N__19718),
            .in3(N__19709),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__19706),
            .in2(N__19691),
            .in3(N__19682),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__19679),
            .in2(N__19664),
            .in3(N__19655),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__19652),
            .in2(N__19637),
            .in3(N__19628),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__19625),
            .in2(N__19613),
            .in3(N__19598),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__19595),
            .in2(N__19589),
            .in3(N__19571),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__19787),
            .in2(N__19568),
            .in3(N__19550),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__19790),
            .in2(N__19547),
            .in3(N__19529),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__19788),
            .in2(N__19865),
            .in3(N__19847),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__19791),
            .in2(N__19844),
            .in3(N__19826),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__19789),
            .in2(N__19823),
            .in3(N__19805),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__19792),
            .in2(N__19763),
            .in3(N__19751),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_15_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_15_0  (
            .in0(N__19748),
            .in1(N__20864),
            .in2(_gnd_net_),
            .in3(N__19736),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_1_15_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_1_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_1_15_1  (
            .in0(N__20085),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20641),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_1_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_1_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27628),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3  (
            .in0(N__20128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20665),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_5  (
            .in0(N__20161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20695),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_1_15_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_1_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_1_15_7  (
            .in0(N__20362),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20611),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_16_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_16_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__19882),
            .in2(_gnd_net_),
            .in3(N__20203),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_1_16_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_1_16_1 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_1_16_1  (
            .in0(N__19883),
            .in1(N__21195),
            .in2(N__19868),
            .in3(N__20189),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_1_16_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_1_16_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_1_16_2  (
            .in0(N__20702),
            .in1(N__20141),
            .in2(N__21219),
            .in3(N__20160),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_1_16_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_1_16_3 .LUT_INIT=16'b1011100001110100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_1_16_3  (
            .in0(N__21125),
            .in1(N__21196),
            .in2(N__21146),
            .in3(N__20174),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_1_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_1_16_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_1_16_4  (
            .in0(N__20669),
            .in1(N__20108),
            .in2(N__21220),
            .in3(N__20127),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_1_16_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_1_16_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_1_16_5  (
            .in0(N__20615),
            .in1(N__21204),
            .in2(N__20342),
            .in3(N__20361),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_1_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_1_16_6 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_1_16_6  (
            .in0(N__21203),
            .in1(N__20645),
            .in2(N__20089),
            .in3(N__20063),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_1_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_1_16_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_1_16_7  (
            .in0(N__21062),
            .in1(N__20327),
            .in2(N__21230),
            .in3(N__21044),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_1_18_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_1_18_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_1_18_4  (
            .in0(N__21104),
            .in1(N__21218),
            .in2(N__21086),
            .in3(N__20315),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_19_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__20036),
            .in2(_gnd_net_),
            .in3(N__20051),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_19_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__20018),
            .in2(_gnd_net_),
            .in3(N__20030),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_19_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__19997),
            .in2(_gnd_net_),
            .in3(N__20012),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_19_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(N__19973),
            .in2(_gnd_net_),
            .in3(N__19991),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_19_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_19_4  (
            .in0(_gnd_net_),
            .in1(N__19952),
            .in2(_gnd_net_),
            .in3(N__19967),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_19_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(N__19931),
            .in2(_gnd_net_),
            .in3(N__19946),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_19_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(N__19910),
            .in2(_gnd_net_),
            .in3(N__19925),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_19_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__19889),
            .in2(_gnd_net_),
            .in3(N__19904),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_20_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(N__20231),
            .in2(_gnd_net_),
            .in3(N__20246),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_20_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(N__20213),
            .in2(_gnd_net_),
            .in3(N__20225),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_20_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_20_2  (
            .in0(_gnd_net_),
            .in1(N__20207),
            .in2(_gnd_net_),
            .in3(N__20180),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_1_20_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_1_20_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_1_20_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_1_20_3  (
            .in0(N__21214),
            .in1(N__20756),
            .in2(_gnd_net_),
            .in3(N__20177),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_20_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(N__21120),
            .in2(_gnd_net_),
            .in3(N__20165),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_20_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_20_5  (
            .in0(_gnd_net_),
            .in1(N__20162),
            .in2(_gnd_net_),
            .in3(N__20132),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_20_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_20_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_20_6  (
            .in0(_gnd_net_),
            .in1(N__20129),
            .in2(_gnd_net_),
            .in3(N__20093),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_20_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20090),
            .in3(N__20054),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_21_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_21_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_21_0  (
            .in0(_gnd_net_),
            .in1(N__20366),
            .in2(_gnd_net_),
            .in3(N__20330),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_21_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_21_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_21_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_21_1  (
            .in0(_gnd_net_),
            .in1(N__21036),
            .in2(_gnd_net_),
            .in3(N__20318),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_21_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_21_2  (
            .in0(_gnd_net_),
            .in1(N__21081),
            .in2(_gnd_net_),
            .in3(N__20306),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_21_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_21_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20303),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.N_42_i_i_LC_1_30_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.N_42_i_i_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.N_42_i_i_LC_1_30_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst1.N_42_i_i_LC_1_30_1  (
            .in0(_gnd_net_),
            .in1(N__35066),
            .in2(_gnd_net_),
            .in3(N__48682),
            .lcout(N_42_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2  (
            .in0(N__20521),
            .in1(N__20494),
            .in2(N__20272),
            .in3(N__20294),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_2_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_2_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_2_10_4 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_2_10_4  (
            .in0(N__23188),
            .in1(N__22296),
            .in2(N__22619),
            .in3(N__22409),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49145),
            .ce(),
            .sr(N__48630));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_11_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_11_0  (
            .in0(N__20566),
            .in1(N__20583),
            .in2(N__20548),
            .in3(N__20288),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_11_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_11_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__20287),
            .in2(_gnd_net_),
            .in3(N__20265),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_11_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_11_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_11_3  (
            .in0(N__20584),
            .in1(N__20567),
            .in2(N__20552),
            .in3(N__20544),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_11_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_11_4 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_2_11_4  (
            .in0(N__20432),
            .in1(N__20520),
            .in2(N__20501),
            .in3(N__20493),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_11_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_11_6  (
            .in0(N__20470),
            .in1(N__20456),
            .in2(_gnd_net_),
            .in3(N__20444),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_12_3 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_12_3  (
            .in0(N__20770),
            .in1(N__23168),
            .in2(N__22712),
            .in3(N__22280),
            .lcout(\current_shift_inst.PI_CTRL.N_140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_6 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_6  (
            .in0(N__23167),
            .in1(N__22707),
            .in2(_gnd_net_),
            .in3(N__20769),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_7 .LUT_INIT=16'b0101010100010000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_7  (
            .in0(N__22753),
            .in1(N__22281),
            .in2(N__20408),
            .in3(N__21453),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_13_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_13_1  (
            .in0(N__23169),
            .in1(N__20771),
            .in2(_gnd_net_),
            .in3(N__22279),
            .lcout(\current_shift_inst.PI_CTRL.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__22956),
            .in2(_gnd_net_),
            .in3(N__22654),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_13_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_13_7  (
            .in0(N__22564),
            .in1(N__22612),
            .in2(N__20774),
            .in3(N__22538),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__20752),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__20729),
            .in2(_gnd_net_),
            .in3(N__20717),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__20714),
            .in2(_gnd_net_),
            .in3(N__20684),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__20681),
            .in2(_gnd_net_),
            .in3(N__20654),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__20651),
            .in2(_gnd_net_),
            .in3(N__20630),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__44868),
            .in2(N__20627),
            .in3(N__20600),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__20597),
            .in2(N__44924),
            .in3(N__20591),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__44872),
            .in2(N__20852),
            .in3(N__20840),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__20837),
            .in2(_gnd_net_),
            .in3(N__20828),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__20825),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__20816),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__20807),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__20798),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__20792),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__20786),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__20780),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__20903),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__20894),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__20885),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__20876),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20867),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_2_16_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_2_16_5 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_2_16_5  (
            .in0(N__22109),
            .in1(N__20987),
            .in2(N__22057),
            .in3(N__21881),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_2_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_2_16_6 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_2_16_6  (
            .in0(N__21882),
            .in1(N__22040),
            .in2(N__22118),
            .in3(N__20972),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_2_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_2_16_7 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_2_16_7  (
            .in0(N__22110),
            .in1(N__20939),
            .in2(N__22058),
            .in3(N__21883),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_2_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_2_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__20858),
            .in2(N__21238),
            .in3(N__21234),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31 ),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_2_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_2_17_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20999),
            .in3(N__20981),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_2_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_2_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__20978),
            .in2(_gnd_net_),
            .in3(N__20966),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_2_17_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_2_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__20963),
            .in2(_gnd_net_),
            .in3(N__20957),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_2_17_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_2_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__20954),
            .in2(_gnd_net_),
            .in3(N__20948),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_2_17_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_2_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__20945),
            .in2(_gnd_net_),
            .in3(N__20933),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_2_17_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_2_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__20930),
            .in2(_gnd_net_),
            .in3(N__20924),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_2_17_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_2_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__20921),
            .in2(_gnd_net_),
            .in3(N__20915),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_2_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_2_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_2_18_0  (
            .in0(_gnd_net_),
            .in1(N__20912),
            .in2(_gnd_net_),
            .in3(N__20906),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271 ),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_2_18_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_2_18_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_2_18_1  (
            .in0(N__21257),
            .in1(N__21248),
            .in2(N__21239),
            .in3(N__21149),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_19_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_19_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__21139),
            .in2(_gnd_net_),
            .in3(N__21124),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_20_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_20_0  (
            .in0(_gnd_net_),
            .in1(N__21082),
            .in2(_gnd_net_),
            .in3(N__21100),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_20_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_20_4  (
            .in0(N__21040),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21061),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_2_30_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_2_30_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_2_30_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \phase_controller_inst1.un7_start_stop_0_a2_LC_2_30_1  (
            .in0(_gnd_net_),
            .in1(N__35065),
            .in2(_gnd_net_),
            .in3(N__48681),
            .lcout(un7_start_stop_0_a2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_3_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_3_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_3_9_3  (
            .in0(_gnd_net_),
            .in1(N__21283),
            .in2(_gnd_net_),
            .in3(N__21379),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_3_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_3_9_4 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_3_9_4  (
            .in0(N__21757),
            .in1(N__21799),
            .in2(N__21011),
            .in3(N__21331),
            .lcout(\pwm_generator_inst.un1_counterlt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_3_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_3_10_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_3_10_3  (
            .in0(N__21550),
            .in1(N__21582),
            .in2(_gnd_net_),
            .in3(N__21628),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto9_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_3_10_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_3_10_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_3_10_4  (
            .in0(N__21665),
            .in1(N__21715),
            .in2(N__21008),
            .in3(N__21005),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_13_7 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_13_7  (
            .in0(N__23166),
            .in1(N__21814),
            .in2(N__21419),
            .in3(N__22376),
            .lcout(\current_shift_inst.PI_CTRL.N_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_3_14_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_3_14_2 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_3_14_2  (
            .in0(N__21863),
            .in1(N__22099),
            .in2(N__22061),
            .in3(N__21437),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_3_14_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_3_14_5 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_3_14_5  (
            .in0(N__22097),
            .in1(N__21428),
            .in2(N__22060),
            .in3(N__21862),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(N__22703),
            .in2(_gnd_net_),
            .in3(N__22752),
            .lcout(\current_shift_inst.PI_CTRL.N_146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_3_14_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_3_14_7 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_3_14_7  (
            .in0(N__22098),
            .in1(N__22053),
            .in2(N__21410),
            .in3(N__21864),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__21353),
            .in2(N__21395),
            .in3(N__21383),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__21305),
            .in2(N__21347),
            .in3(N__21335),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__21263),
            .in2(N__21299),
            .in3(N__21290),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__21776),
            .in2(N__21839),
            .in3(N__21803),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__21731),
            .in2(N__21770),
            .in3(N__21761),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__21683),
            .in2(N__21725),
            .in3(N__21716),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__21635),
            .in2(N__21677),
            .in3(N__21664),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__21596),
            .in2(N__22130),
            .in3(N__21629),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__21563),
            .in2(N__22145),
            .in3(N__21590),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(N__21530),
            .in2(N__22163),
            .in3(N__21557),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_3_16_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_3_16_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_3_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21524),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49109),
            .ce(),
            .sr(N__48652));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_3_17_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_3_17_0 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_3_17_0  (
            .in0(N__22117),
            .in1(N__21887),
            .in2(N__22172),
            .in3(N__22049),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_3_17_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_3_17_2 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_3_17_2  (
            .in0(N__22116),
            .in1(N__22048),
            .in2(N__22154),
            .in3(N__21886),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_3_17_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_3_17_3 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_3_17_3  (
            .in0(N__21885),
            .in1(N__22115),
            .in2(N__22059),
            .in3(N__22136),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_3_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_3_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27422),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_17_6 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_17_6  (
            .in0(N__22114),
            .in1(N__22044),
            .in2(N__21896),
            .in3(N__21884),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_13_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_13_3  (
            .in0(N__22530),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22647),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_13_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_13_4  (
            .in0(N__22605),
            .in1(N__22563),
            .in2(N__21827),
            .in3(N__22957),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_4_13_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_13_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_13_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_14_2  (
            .in0(N__22487),
            .in1(N__22430),
            .in2(N__22343),
            .in3(N__22328),
            .lcout(\current_shift_inst.PI_CTRL.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_4_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_4_14_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_4_14_7  (
            .in0(N__28301),
            .in1(N__30095),
            .in2(N__27430),
            .in3(N__32032),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_4_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_4_15_0 .LUT_INIT=16'b1111111100001011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_4_15_0  (
            .in0(N__22202),
            .in1(N__25018),
            .in2(N__27206),
            .in3(N__22208),
            .lcout(\current_shift_inst.PI_CTRL.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_4_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_4_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_4_15_2  (
            .in0(N__29766),
            .in1(N__27813),
            .in2(N__29834),
            .in3(N__29914),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_4_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_4_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_4_15_3  (
            .in0(N__22226),
            .in1(N__22445),
            .in2(N__22220),
            .in3(N__22217),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_4_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_4_15_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__24205),
            .in2(_gnd_net_),
            .in3(N__27153),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_4_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_4_15_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_4_15_5  (
            .in0(N__27862),
            .in1(N__31856),
            .in2(N__22211),
            .in3(N__27529),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_4_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_4_15_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_4_15_7  (
            .in0(N__27259),
            .in1(N__27104),
            .in2(_gnd_net_),
            .in3(N__26959),
            .lcout(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__22885),
            .in2(_gnd_net_),
            .in3(N__22921),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_16_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_16_1  (
            .in0(N__22993),
            .in1(N__23006),
            .in2(N__23237),
            .in3(N__23038),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_16_2  (
            .in0(N__23258),
            .in1(N__22909),
            .in2(N__22421),
            .in3(N__22418),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_16_3  (
            .in0(N__22310),
            .in1(N__22349),
            .in2(N__22412),
            .in3(N__22316),
            .lcout(\current_shift_inst.PI_CTRL.N_164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_16_4  (
            .in0(N__23071),
            .in1(N__22849),
            .in2(N__23057),
            .in3(N__22861),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_5  (
            .in0(N__22862),
            .in1(N__22850),
            .in2(N__22994),
            .in3(N__23005),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6  (
            .in0(N__23233),
            .in1(N__22922),
            .in2(N__22820),
            .in3(N__22835),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7  (
            .in0(N__22910),
            .in1(N__22889),
            .in2(N__22331),
            .in3(N__22454),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_17_0  (
            .in0(_gnd_net_),
            .in1(N__22816),
            .in2(_gnd_net_),
            .in3(N__22834),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_17_1  (
            .in0(N__23024),
            .in1(N__22975),
            .in2(N__22319),
            .in3(N__23287),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_17_2  (
            .in0(N__23272),
            .in1(N__23111),
            .in2(N__23099),
            .in3(N__23216),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_3  (
            .in0(N__23110),
            .in1(_gnd_net_),
            .in2(N__23095),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_4_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_4_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27692),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_4_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_4_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_4_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_4_17_6  (
            .in0(N__27371),
            .in1(N__27693),
            .in2(N__41284),
            .in3(N__27744),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_4_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_4_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_4_17_7  (
            .in0(N__24140),
            .in1(N__24149),
            .in2(N__22448),
            .in3(N__24167),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_4_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_4_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_4_18_1  (
            .in0(_gnd_net_),
            .in1(N__28293),
            .in2(_gnd_net_),
            .in3(N__27423),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_4_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_4_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_4_18_2  (
            .in0(N__22493),
            .in1(N__25498),
            .in2(N__22436),
            .in3(N__30089),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(N__23215),
            .in2(_gnd_net_),
            .in3(N__23273),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_18_4  (
            .in0(N__23251),
            .in1(N__23020),
            .in2(N__22433),
            .in3(N__23039),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_4_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_4_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_4_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27365),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_4_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_4_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_4_18_6  (
            .in0(N__29910),
            .in1(N__29756),
            .in2(N__29835),
            .in3(N__27809),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_18_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_18_7  (
            .in0(N__23056),
            .in1(N__22976),
            .in2(N__23075),
            .in3(N__23288),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_5_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_5_9_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__26795),
            .in2(_gnd_net_),
            .in3(N__24722),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_5_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_5_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_5_9_2 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_5_9_2  (
            .in0(N__26743),
            .in1(N__24695),
            .in2(N__22478),
            .in3(N__23532),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49138),
            .ce(),
            .sr(N__48598));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_5_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_5_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_5_10_2  (
            .in0(N__26826),
            .in1(N__28558),
            .in2(_gnd_net_),
            .in3(N__34608),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_5_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_5_11_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_5_11_0  (
            .in0(N__23893),
            .in1(N__22475),
            .in2(N__24131),
            .in3(N__22463),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_5_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_5_11_1 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_5_11_1  (
            .in0(N__22462),
            .in1(N__22474),
            .in2(N__23897),
            .in3(N__24130),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_5_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_5_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_29_LC_5_12_0  (
            .in0(N__26827),
            .in1(N__28562),
            .in2(_gnd_net_),
            .in3(N__34686),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49125),
            .ce(N__24806),
            .sr(N__48623));
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_5_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_5_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_28_LC_5_12_7  (
            .in0(N__34685),
            .in1(N__26876),
            .in2(_gnd_net_),
            .in3(N__26894),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49125),
            .ce(N__24806),
            .sr(N__48623));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33922),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49119),
            .ce(),
            .sr(N__48631));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33092),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48637));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33388),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48637));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33842),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48637));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33298),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48637));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33056),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48637));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_5  (
            .in0(N__33186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48637));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33011),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48637));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33887),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48637));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__23960),
            .in2(N__26960),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__49102),
            .ce(),
            .sr(N__48640));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__22802),
            .in2(N__27103),
            .in3(N__22784),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__49102),
            .ce(),
            .sr(N__48640));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__22781),
            .in2(N__27260),
            .in3(N__22763),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__49102),
            .ce(),
            .sr(N__48640));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__33137),
            .in2(N__25019),
            .in3(N__22724),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__49102),
            .ce(),
            .sr(N__48640));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__27202),
            .in2(N__22721),
            .in3(N__22670),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__49102),
            .ce(),
            .sr(N__48640));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_5  (
            .in0(_gnd_net_),
            .in1(N__22667),
            .in2(N__27158),
            .in3(N__22628),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__49102),
            .ce(),
            .sr(N__48640));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(N__22625),
            .in2(N__27866),
            .in3(N__22580),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__49102),
            .ce(),
            .sr(N__48640));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(N__22577),
            .in2(N__24209),
            .in3(N__22541),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__49102),
            .ce(),
            .sr(N__48640));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(N__33749),
            .in2(N__27530),
            .in3(N__22508),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__49094),
            .ce(),
            .sr(N__48644));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(N__31814),
            .in2(N__31868),
            .in3(N__22934),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__49094),
            .ce(),
            .sr(N__48644));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(N__22931),
            .in2(N__28235),
            .in3(N__22913),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__49094),
            .ce(),
            .sr(N__48644));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(N__41283),
            .in2(N__23123),
            .in3(N__22901),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__49094),
            .ce(),
            .sr(N__48644));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(N__22898),
            .in2(N__27431),
            .in3(N__22874),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__49094),
            .ce(),
            .sr(N__48644));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_5  (
            .in0(_gnd_net_),
            .in1(N__22871),
            .in2(N__29915),
            .in3(N__22853),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__49094),
            .ce(),
            .sr(N__48644));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(N__31778),
            .in2(N__27817),
            .in3(N__22838),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__49094),
            .ce(),
            .sr(N__48644));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(N__27695),
            .in2(N__31796),
            .in3(N__22823),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__49094),
            .ce(),
            .sr(N__48644));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(N__31733),
            .in2(N__29840),
            .in3(N__22805),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_5_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__49085),
            .ce(),
            .sr(N__48648));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(N__27370),
            .in2(N__31757),
            .in3(N__23102),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__49085),
            .ce(),
            .sr(N__48648));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(N__31737),
            .in2(N__27638),
            .in3(N__23078),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__49085),
            .ce(),
            .sr(N__48648));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(N__35471),
            .in2(N__31758),
            .in3(N__23060),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__49085),
            .ce(),
            .sr(N__48648));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(N__31741),
            .in2(N__27749),
            .in3(N__23042),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__49085),
            .ce(),
            .sr(N__48648));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(N__27574),
            .in2(N__31759),
            .in3(N__23027),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__49085),
            .ce(),
            .sr(N__48648));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_6  (
            .in0(_gnd_net_),
            .in1(N__31745),
            .in2(N__29984),
            .in3(N__23009),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__49085),
            .ce(),
            .sr(N__48648));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(N__29767),
            .in2(N__31760),
            .in3(N__22997),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__49085),
            .ce(),
            .sr(N__48648));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(N__31782),
            .in2(N__28064),
            .in3(N__22979),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_5_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__49077),
            .ce(),
            .sr(N__48653));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(N__28012),
            .in2(N__31797),
            .in3(N__22964),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__49077),
            .ce(),
            .sr(N__48653));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__31786),
            .in2(N__27950),
            .in3(N__23276),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__49077),
            .ce(),
            .sr(N__48653));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(N__30090),
            .in2(N__31798),
            .in3(N__23261),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__49077),
            .ce(),
            .sr(N__48653));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(N__31790),
            .in2(N__25502),
            .in3(N__23240),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__49077),
            .ce(),
            .sr(N__48653));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(N__42757),
            .in2(N__31799),
            .in3(N__23219),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__49077),
            .ce(),
            .sr(N__48653));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(N__31794),
            .in2(N__28297),
            .in3(N__23204),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__49077),
            .ce(),
            .sr(N__48653));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_7  (
            .in0(N__31795),
            .in1(N__32033),
            .in2(_gnd_net_),
            .in3(N__23201),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49077),
            .ce(),
            .sr(N__48653));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33523),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49070),
            .ce(),
            .sr(N__48657));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_7_0  (
            .in0(N__34484),
            .in1(N__30403),
            .in2(_gnd_net_),
            .in3(N__30382),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_7_3  (
            .in0(N__30151),
            .in1(N__30130),
            .in2(_gnd_net_),
            .in3(N__34483),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_7_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_7_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_7_7_5  (
            .in0(N__32731),
            .in1(N__32707),
            .in2(_gnd_net_),
            .in3(N__34482),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_8_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_8_0  (
            .in0(N__23767),
            .in1(N__23743),
            .in2(N__23300),
            .in3(N__23309),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_7_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_7_8_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_7_8_1  (
            .in0(N__23308),
            .in1(N__23768),
            .in2(N__23747),
            .in3(N__23296),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_7_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_7_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_7_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_7_8_2  (
            .in0(N__28952),
            .in1(N__28973),
            .in2(_gnd_net_),
            .in3(N__34693),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49134),
            .ce(N__24801),
            .sr(N__48570));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_7_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_7_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_7_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_7_8_3  (
            .in0(N__34688),
            .in1(N__29012),
            .in2(_gnd_net_),
            .in3(N__29033),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49134),
            .ce(N__24801),
            .sr(N__48570));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_7_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_7_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_7_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_7_8_4  (
            .in0(N__29188),
            .in1(N__29205),
            .in2(_gnd_net_),
            .in3(N__34694),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49134),
            .ce(N__24801),
            .sr(N__48570));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_7_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_7_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_7_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_7_8_5  (
            .in0(N__34689),
            .in1(N__30274),
            .in2(_gnd_net_),
            .in3(N__30242),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49134),
            .ce(N__24801),
            .sr(N__48570));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_7_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_7_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_7_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_7_8_6  (
            .in0(N__28463),
            .in1(N__28433),
            .in2(_gnd_net_),
            .in3(N__34695),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49134),
            .ce(N__24801),
            .sr(N__48570));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_7_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_7_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_7_8_7 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_7_8_7  (
            .in0(N__30147),
            .in1(N__30126),
            .in2(N__34706),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49134),
            .ce(N__24801),
            .sr(N__48570));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_7_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_7_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__24533),
            .in2(N__23417),
            .in3(N__23533),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_7_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_7_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__24527),
            .in2(N__23408),
            .in3(N__23513),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_7_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_7_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__24521),
            .in2(N__23399),
            .in3(N__23720),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_7_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_7_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(N__23390),
            .in2(N__23381),
            .in3(N__23702),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_7_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_7_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__23372),
            .in2(N__23366),
            .in3(N__23684),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_7_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_7_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_7_9_5  (
            .in0(N__23663),
            .in1(N__23357),
            .in2(N__23348),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_7_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_7_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__23336),
            .in2(N__23330),
            .in3(N__23642),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_7_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_7_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(N__24425),
            .in2(N__23321),
            .in3(N__23624),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_7_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_7_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__24407),
            .in2(N__23495),
            .in3(N__23606),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_7_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_7_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__23486),
            .in2(N__24398),
            .in3(N__23585),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_7_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_7_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__23480),
            .in2(N__24551),
            .in3(N__23867),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_7_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_7_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(N__24557),
            .in2(N__23474),
            .in3(N__23849),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_7_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_7_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__24440),
            .in2(N__23465),
            .in3(N__23831),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_7_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_7_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_7_10_5  (
            .in0(N__23810),
            .in1(N__24647),
            .in2(N__23456),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_7_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_7_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__23444),
            .in2(N__24542),
            .in3(N__23792),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_7_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_7_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__24329),
            .in2(N__24386),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_7_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_7_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__23438),
            .in2(N__23429),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_7_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_7_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__24239),
            .in2(N__24299),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_7_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_7_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__24587),
            .in2(N__24641),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_7_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_7_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__24974),
            .in2(N__24917),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_7_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_7_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__24902),
            .in2(N__24845),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_7_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_7_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__23564),
            .in2(N__23555),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_7_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_7_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__24754),
            .in2(N__24452),
            .in3(N__23543),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_7_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_7_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23540),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__23537),
            .in2(N__24731),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_12_1  (
            .in0(N__24046),
            .in1(N__23512),
            .in2(_gnd_net_),
            .in3(N__23498),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49111),
            .ce(),
            .sr(N__48606));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_12_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_12_2  (
            .in0(N__24050),
            .in1(N__23719),
            .in2(N__24677),
            .in3(N__23705),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49111),
            .ce(),
            .sr(N__48606));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_12_3  (
            .in0(N__24047),
            .in1(N__23701),
            .in2(_gnd_net_),
            .in3(N__23687),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49111),
            .ce(),
            .sr(N__48606));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_12_4  (
            .in0(N__24051),
            .in1(N__23680),
            .in2(_gnd_net_),
            .in3(N__23666),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49111),
            .ce(),
            .sr(N__48606));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_12_5  (
            .in0(N__24048),
            .in1(N__23659),
            .in2(_gnd_net_),
            .in3(N__23645),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49111),
            .ce(),
            .sr(N__48606));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_12_6  (
            .in0(N__24052),
            .in1(N__23641),
            .in2(_gnd_net_),
            .in3(N__23627),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49111),
            .ce(),
            .sr(N__48606));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_12_7  (
            .in0(N__24049),
            .in1(N__23623),
            .in2(_gnd_net_),
            .in3(N__23609),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49111),
            .ce(),
            .sr(N__48606));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_13_0  (
            .in0(N__24045),
            .in1(N__23602),
            .in2(_gnd_net_),
            .in3(N__23588),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49103),
            .ce(),
            .sr(N__48616));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_13_1  (
            .in0(N__24038),
            .in1(N__23581),
            .in2(_gnd_net_),
            .in3(N__23567),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49103),
            .ce(),
            .sr(N__48616));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_13_2  (
            .in0(N__24042),
            .in1(N__23866),
            .in2(_gnd_net_),
            .in3(N__23852),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49103),
            .ce(),
            .sr(N__48616));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_13_3  (
            .in0(N__24039),
            .in1(N__23848),
            .in2(_gnd_net_),
            .in3(N__23834),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49103),
            .ce(),
            .sr(N__48616));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_13_4  (
            .in0(N__24043),
            .in1(N__23827),
            .in2(_gnd_net_),
            .in3(N__23813),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49103),
            .ce(),
            .sr(N__48616));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_13_5  (
            .in0(N__24040),
            .in1(N__23809),
            .in2(_gnd_net_),
            .in3(N__23795),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49103),
            .ce(),
            .sr(N__48616));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_13_6  (
            .in0(N__24044),
            .in1(N__23791),
            .in2(_gnd_net_),
            .in3(N__23777),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49103),
            .ce(),
            .sr(N__48616));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_13_7  (
            .in0(N__24041),
            .in1(N__24370),
            .in2(_gnd_net_),
            .in3(N__23774),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49103),
            .ce(),
            .sr(N__48616));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_14_0  (
            .in0(N__24087),
            .in1(N__24343),
            .in2(_gnd_net_),
            .in3(N__23771),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49095),
            .ce(),
            .sr(N__48624));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_14_1  (
            .in0(N__24098),
            .in1(N__23766),
            .in2(_gnd_net_),
            .in3(N__23750),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49095),
            .ce(),
            .sr(N__48624));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_14_2  (
            .in0(N__24088),
            .in1(N__23737),
            .in2(_gnd_net_),
            .in3(N__23723),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49095),
            .ce(),
            .sr(N__48624));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_14_3  (
            .in0(N__24099),
            .in1(N__24277),
            .in2(_gnd_net_),
            .in3(N__23921),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49095),
            .ce(),
            .sr(N__48624));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_14_4  (
            .in0(N__24089),
            .in1(N__24253),
            .in2(_gnd_net_),
            .in3(N__23918),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49095),
            .ce(),
            .sr(N__48624));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_14_5  (
            .in0(N__24100),
            .in1(N__24627),
            .in2(_gnd_net_),
            .in3(N__23915),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49095),
            .ce(),
            .sr(N__48624));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_14_6  (
            .in0(N__24090),
            .in1(N__24601),
            .in2(_gnd_net_),
            .in3(N__23912),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49095),
            .ce(),
            .sr(N__48624));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_14_7  (
            .in0(N__24101),
            .in1(N__24953),
            .in2(_gnd_net_),
            .in3(N__23909),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49095),
            .ce(),
            .sr(N__48624));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_15_0  (
            .in0(N__24091),
            .in1(N__24933),
            .in2(_gnd_net_),
            .in3(N__23906),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49086),
            .ce(),
            .sr(N__48632));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_15_1  (
            .in0(N__24095),
            .in1(N__24891),
            .in2(_gnd_net_),
            .in3(N__23903),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49086),
            .ce(),
            .sr(N__48632));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_15_2  (
            .in0(N__24092),
            .in1(N__24870),
            .in2(_gnd_net_),
            .in3(N__23900),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49086),
            .ce(),
            .sr(N__48632));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_15_3  (
            .in0(N__24096),
            .in1(N__23886),
            .in2(_gnd_net_),
            .in3(N__23870),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49086),
            .ce(),
            .sr(N__48632));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_15_4  (
            .in0(N__24093),
            .in1(N__24121),
            .in2(_gnd_net_),
            .in3(N__24107),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49086),
            .ce(),
            .sr(N__48632));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_15_5  (
            .in0(N__24097),
            .in1(N__24466),
            .in2(_gnd_net_),
            .in3(N__24104),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49086),
            .ce(),
            .sr(N__48632));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_15_6  (
            .in0(N__24094),
            .in1(N__24490),
            .in2(_gnd_net_),
            .in3(N__23963),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49086),
            .ce(),
            .sr(N__48632));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_7_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_7_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_7_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33722),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49086),
            .ce(),
            .sr(N__48632));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_7_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_7_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_7_16_0  (
            .in0(N__24173),
            .in1(N__23951),
            .in2(N__24158),
            .in3(N__23933),
            .lcout(\current_shift_inst.PI_CTRL.N_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_16_2  (
            .in0(N__27518),
            .in1(N__27861),
            .in2(N__31864),
            .in3(N__24204),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_16_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_16_3  (
            .in0(N__27200),
            .in1(N__25008),
            .in2(N__23939),
            .in3(N__27149),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_72_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_7_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_7_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_7_16_4  (
            .in0(N__23927),
            .in1(N__42753),
            .in2(N__23936),
            .in3(N__28233),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_7_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_7_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_7_16_5  (
            .in0(N__27685),
            .in1(N__41266),
            .in2(N__27369),
            .in3(N__27743),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_7_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_7_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_7_17_0  (
            .in0(N__29966),
            .in1(N__27630),
            .in2(N__35474),
            .in3(N__32009),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_17_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__42749),
            .in2(_gnd_net_),
            .in3(N__28229),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_7_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_7_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28292),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_17_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_17_3  (
            .in0(N__27939),
            .in1(N__28004),
            .in2(N__28060),
            .in3(N__27560),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_7_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_7_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_7_17_4  (
            .in0(N__29965),
            .in1(N__27629),
            .in2(N__35473),
            .in3(N__28053),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30076),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_7_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_7_17_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_7_17_7  (
            .in0(N__27938),
            .in1(N__25491),
            .in2(N__28011),
            .in3(N__27559),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_7_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_7_18_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_7_18_0  (
            .in0(N__24189),
            .in1(N__33524),
            .in2(N__35405),
            .in3(N__29486),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_7_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_7_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24188),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_7_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_7_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_7_18_2 .LUT_INIT=16'b0000111100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_7_18_2  (
            .in0(N__32199),
            .in1(N__32022),
            .in2(N__25139),
            .in3(N__32381),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49065),
            .ce(),
            .sr(N__48645));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_7_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_7_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_7_18_3 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_7_18_3  (
            .in0(N__32018),
            .in1(N__32200),
            .in2(N__32398),
            .in3(N__25211),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49065),
            .ce(),
            .sr(N__48645));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_7_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_7_18_4 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_7_18_4  (
            .in0(N__32197),
            .in1(N__32020),
            .in2(N__25436),
            .in3(N__32379),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49065),
            .ce(),
            .sr(N__48645));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_7_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_7_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_7_18_5 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_7_18_5  (
            .in0(N__32019),
            .in1(N__32201),
            .in2(N__32399),
            .in3(N__25424),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49065),
            .ce(),
            .sr(N__48645));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_18_6 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_7_18_6  (
            .in0(N__32198),
            .in1(N__32021),
            .in2(N__25415),
            .in3(N__32380),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49065),
            .ce(),
            .sr(N__48645));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27131),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_7_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_7_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_7_19_2 .LUT_INIT=16'b0000111100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_7_19_2  (
            .in0(N__32192),
            .in1(N__32004),
            .in2(N__25175),
            .in3(N__32365),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49059),
            .ce(),
            .sr(N__48649));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_19_5 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_7_19_5  (
            .in0(N__32003),
            .in1(N__32193),
            .in2(N__32396),
            .in3(N__25367),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49059),
            .ce(),
            .sr(N__48649));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_7_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_7_19_6 .LUT_INIT=16'b0100010001010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_7_19_6  (
            .in0(N__25118),
            .in1(N__32366),
            .in2(N__32219),
            .in3(N__32005),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49059),
            .ce(),
            .sr(N__48649));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_7_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_7_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27499),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_7_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_7_20_2 .LUT_INIT=16'b0010001011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_7_20_2  (
            .in0(N__32028),
            .in1(N__32369),
            .in2(N__32223),
            .in3(N__25358),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49051),
            .ce(),
            .sr(N__48654));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_7_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_7_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_7_20_3 .LUT_INIT=16'b0100111101001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_7_20_3  (
            .in0(N__32367),
            .in1(N__32029),
            .in2(N__25400),
            .in3(N__32211),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49051),
            .ce(),
            .sr(N__48654));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_20_5 .LUT_INIT=16'b0100111101001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_7_20_5  (
            .in0(N__32368),
            .in1(N__32030),
            .in2(N__25388),
            .in3(N__32212),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49051),
            .ce(),
            .sr(N__48654));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_7_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_7_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_7_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27733),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_8_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_8_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_8_5_5 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_8_5_5  (
            .in0(N__24227),
            .in1(N__28154),
            .in2(_gnd_net_),
            .in3(N__28187),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49142),
            .ce(),
            .sr(N__48537));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_8_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_8_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24224),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_6_3  (
            .in0(N__34609),
            .in1(N__28462),
            .in2(_gnd_net_),
            .in3(N__28422),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_8_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_8_6_4 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__24226),
            .in2(N__28186),
            .in3(N__28150),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_204_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_6_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_6_7  (
            .in0(N__24225),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28179),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_203_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_7_0  (
            .in0(N__29234),
            .in1(N__29288),
            .in2(N__29184),
            .in3(N__28814),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_7_1 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__26875),
            .in2(N__24302),
            .in3(N__26431),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25786),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49135),
            .ce(N__26479),
            .sr(N__48550));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_7_3  (
            .in0(N__25760),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49135),
            .ce(N__26479),
            .sr(N__48550));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_7_4  (
            .in0(N__28851),
            .in1(N__28815),
            .in2(_gnd_net_),
            .in3(N__34481),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_8_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_8_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_8_7_5  (
            .in0(N__29289),
            .in1(N__34476),
            .in2(_gnd_net_),
            .in3(N__29325),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_7_6 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_7_6  (
            .in0(N__29235),
            .in1(N__29265),
            .in2(N__34607),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_7_7  (
            .in0(N__34480),
            .in1(N__29209),
            .in2(_gnd_net_),
            .in3(N__29177),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_8_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_8_0  (
            .in0(N__24283),
            .in1(N__24259),
            .in2(N__24419),
            .in3(N__24434),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_8_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_8_1  (
            .in0(N__24433),
            .in1(N__24284),
            .in2(N__24263),
            .in3(N__24415),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_8_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_8_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_20_LC_8_8_2  (
            .in0(N__28895),
            .in1(N__28916),
            .in2(_gnd_net_),
            .in3(N__34672),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49131),
            .ce(N__24800),
            .sr(N__48558));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_8_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_8_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_8_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_8_8_4  (
            .in0(N__30399),
            .in1(N__30375),
            .in2(_gnd_net_),
            .in3(N__34673),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49131),
            .ce(N__24800),
            .sr(N__48558));
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_8_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_8_8_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_21_LC_8_8_5  (
            .in0(N__34768),
            .in1(_gnd_net_),
            .in2(N__34705),
            .in3(N__34744),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49131),
            .ce(N__24800),
            .sr(N__48558));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_6  (
            .in0(N__28337),
            .in1(N__28355),
            .in2(_gnd_net_),
            .in3(N__34674),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49131),
            .ce(N__24800),
            .sr(N__48558));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_7  (
            .in0(N__34668),
            .in1(N__32663),
            .in2(_gnd_net_),
            .in3(N__32634),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49131),
            .ce(N__24800),
            .sr(N__48558));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_8_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_8_9_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_8_9_0  (
            .in0(N__24376),
            .in1(N__24352),
            .in2(N__24314),
            .in3(N__24323),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_8_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_8_9_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_8_9_1  (
            .in0(N__24322),
            .in1(N__24377),
            .in2(N__24356),
            .in3(N__24310),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_8_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_8_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_8_9_2  (
            .in0(N__32777),
            .in1(N__32804),
            .in2(_gnd_net_),
            .in3(N__34679),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49126),
            .ce(N__24802),
            .sr(N__48571));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_8_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_8_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_8_9_3  (
            .in0(N__34675),
            .in1(N__32891),
            .in2(_gnd_net_),
            .in3(N__32921),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49126),
            .ce(N__24802),
            .sr(N__48571));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_8_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_8_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_8_9_4  (
            .in0(N__28631),
            .in1(N__28654),
            .in2(_gnd_net_),
            .in3(N__34678),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49126),
            .ce(N__24802),
            .sr(N__48571));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_8_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_8_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_8_9_5  (
            .in0(N__34676),
            .in1(N__28852),
            .in2(_gnd_net_),
            .in3(N__28822),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49126),
            .ce(N__24802),
            .sr(N__48571));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_6  (
            .in0(N__29326),
            .in1(N__29296),
            .in2(_gnd_net_),
            .in3(N__34680),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49126),
            .ce(N__24802),
            .sr(N__48571));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_7  (
            .in0(N__34677),
            .in1(N__29236),
            .in2(_gnd_net_),
            .in3(N__29266),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49126),
            .ce(N__24802),
            .sr(N__48571));
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_8_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_8_10_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_8_10_0  (
            .in0(N__24474),
            .in1(N__24660),
            .in2(N__24503),
            .in3(N__24514),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_8_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_8_10_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_8_10_1  (
            .in0(N__24513),
            .in1(N__24501),
            .in2(N__24664),
            .in3(N__24475),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_8_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_8_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_30_LC_8_10_2  (
            .in0(N__28493),
            .in1(N__28792),
            .in2(_gnd_net_),
            .in3(N__34616),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49120),
            .ce(N__24803),
            .sr(N__48581));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_10_3 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_10_3  (
            .in0(N__24515),
            .in1(N__24502),
            .in2(N__24665),
            .in3(N__24476),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_10_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_10_4  (
            .in0(N__28687),
            .in1(N__34614),
            .in2(_gnd_net_),
            .in3(N__28674),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_8_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_8_10_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_8_10_5  (
            .in0(N__28675),
            .in1(_gnd_net_),
            .in2(N__24443),
            .in3(N__34622),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49120),
            .ce(N__24803),
            .sr(N__48581));
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_8_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_8_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_31_LC_8_10_6  (
            .in0(N__34623),
            .in1(N__28769),
            .in2(_gnd_net_),
            .in3(N__28744),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49120),
            .ce(N__24803),
            .sr(N__48581));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_8_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_8_10_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_8_10_7  (
            .in0(N__34615),
            .in1(N__32842),
            .in2(_gnd_net_),
            .in3(N__32867),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49120),
            .ce(N__24803),
            .sr(N__48581));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_11_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_11_0  (
            .in0(N__24628),
            .in1(N__24607),
            .in2(N__24572),
            .in3(N__24581),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_8_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_8_11_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_8_11_1  (
            .in0(N__24580),
            .in1(N__24629),
            .in2(N__24611),
            .in3(N__24568),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_8_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_8_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_22_LC_8_11_2  (
            .in0(N__32735),
            .in1(N__32699),
            .in2(_gnd_net_),
            .in3(N__34667),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49112),
            .ce(N__24804),
            .sr(N__48588));
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_8_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_8_11_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_23_LC_8_11_3  (
            .in0(N__34664),
            .in1(_gnd_net_),
            .in2(N__30197),
            .in3(N__30218),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49112),
            .ce(N__24804),
            .sr(N__48588));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_11_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_11_4  (
            .in0(N__28606),
            .in1(N__34662),
            .in2(_gnd_net_),
            .in3(N__28573),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(elapsed_time_ns_1_RNIV8OBB_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_8_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_8_11_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_8_11_5  (
            .in0(N__34663),
            .in1(_gnd_net_),
            .in2(N__24560),
            .in3(N__28607),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49112),
            .ce(N__24804),
            .sr(N__48588));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_8_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_8_11_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_8_11_6  (
            .in0(N__28385),
            .in1(N__34666),
            .in2(_gnd_net_),
            .in3(N__28406),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49112),
            .ce(N__24804),
            .sr(N__48588));
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_8_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_8_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_24_LC_8_11_7  (
            .in0(N__34665),
            .in1(N__29073),
            .in2(_gnd_net_),
            .in3(N__29093),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49112),
            .ce(N__24804),
            .sr(N__48588));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_12_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_12_0  (
            .in0(N__27035),
            .in1(N__35743),
            .in2(N__27053),
            .in3(N__26987),
            .lcout(),
            .ltout(\phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_8_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_8_12_1 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_8_12_1  (
            .in0(N__26678),
            .in1(N__24718),
            .in2(N__24779),
            .in3(N__34841),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49104),
            .ce(),
            .sr(N__48599));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_12_2 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_12_2  (
            .in0(N__26785),
            .in1(N__24775),
            .in2(_gnd_net_),
            .in3(N__24713),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_LC_8_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_8_12_3 .LUT_INIT=16'b1000101011111010;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_8_12_3  (
            .in0(N__24776),
            .in1(N__26758),
            .in2(N__26744),
            .in3(N__26787),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49104),
            .ce(),
            .sr(N__48599));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_8_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_8_12_4 .LUT_INIT=16'b1111110101110101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_8_12_4  (
            .in0(N__26786),
            .in1(N__24767),
            .in2(N__24758),
            .in3(N__24740),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_8_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_8_12_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24734),
            .in3(N__26728),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_8_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_8_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_8_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24714),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49104),
            .ce(),
            .sr(N__48599));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_8_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_8_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__26729),
            .in2(_gnd_net_),
            .in3(N__24688),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_13_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_13_0  (
            .in0(N__24951),
            .in1(N__24934),
            .in2(N__24818),
            .in3(N__24965),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_13_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_13_1  (
            .in0(N__24964),
            .in1(N__24952),
            .in2(N__24938),
            .in3(N__24814),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_13_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_13_2  (
            .in0(N__29446),
            .in1(N__29416),
            .in2(_gnd_net_),
            .in3(N__34696),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_8_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_8_13_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_26_LC_8_13_3  (
            .in0(N__34698),
            .in1(_gnd_net_),
            .in2(N__24905),
            .in3(N__29447),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49096),
            .ce(N__24805),
            .sr(N__48607));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_13_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_13_4  (
            .in0(N__24853),
            .in1(N__24893),
            .in2(N__24875),
            .in3(N__24826),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_13_5 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_13_5  (
            .in0(N__24892),
            .in1(N__24871),
            .in2(N__24830),
            .in3(N__24854),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_8_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_8_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_27_LC_8_13_6  (
            .in0(N__26432),
            .in1(N__26444),
            .in2(_gnd_net_),
            .in3(N__34699),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49096),
            .ce(N__24805),
            .sr(N__48607));
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_8_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_8_13_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_25_LC_8_13_7  (
            .in0(N__34697),
            .in1(N__29141),
            .in2(_gnd_net_),
            .in3(N__29156),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49096),
            .ce(N__24805),
            .sr(N__48607));
    defparam \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_8_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_8_14_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_8_14_0  (
            .in0(N__24993),
            .in1(N__33838),
            .in2(N__35380),
            .in3(N__29534),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24992),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_8_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_8_14_2 .LUT_INIT=16'b0000010111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_8_14_2  (
            .in0(N__32158),
            .in1(_gnd_net_),
            .in2(N__32395),
            .in3(N__25031),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49087),
            .ce(),
            .sr(N__48617));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_8_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_8_14_3 .LUT_INIT=16'b0010001011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_8_14_3  (
            .in0(N__32013),
            .in1(N__32350),
            .in2(N__32202),
            .in3(N__25100),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49087),
            .ce(),
            .sr(N__48617));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_4 .LUT_INIT=16'b0000110011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_4  (
            .in0(N__32156),
            .in1(N__32016),
            .in2(N__32393),
            .in3(N__25079),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49087),
            .ce(),
            .sr(N__48617));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_5 .LUT_INIT=16'b0010001011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_5  (
            .in0(N__32014),
            .in1(N__32351),
            .in2(N__32203),
            .in3(N__25349),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49087),
            .ce(),
            .sr(N__48617));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_8_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_8_14_6 .LUT_INIT=16'b0000110011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_8_14_6  (
            .in0(N__32157),
            .in1(N__32017),
            .in2(N__32394),
            .in3(N__25337),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49087),
            .ce(),
            .sr(N__48617));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_7 .LUT_INIT=16'b0010001011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_7  (
            .in0(N__32015),
            .in1(N__32352),
            .in2(N__32204),
            .in3(N__25313),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49087),
            .ce(),
            .sr(N__48617));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_8_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_8_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27193),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_8_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_8_15_2 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_8_15_2  (
            .in0(N__32132),
            .in1(N__32027),
            .in2(N__25196),
            .in3(N__32328),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49078),
            .ce(),
            .sr(N__48625));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_3 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_3  (
            .in0(N__32023),
            .in1(N__32133),
            .in2(N__32382),
            .in3(N__25301),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49078),
            .ce(),
            .sr(N__48625));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_4 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_4  (
            .in0(N__32130),
            .in1(N__32025),
            .in2(N__25280),
            .in3(N__32326),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49078),
            .ce(),
            .sr(N__48625));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_15_5 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_8_15_5  (
            .in0(N__32024),
            .in1(N__32134),
            .in2(N__32383),
            .in3(N__25250),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49078),
            .ce(),
            .sr(N__48625));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_6 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_6  (
            .in0(N__32131),
            .in1(N__32026),
            .in2(N__25238),
            .in3(N__32327),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49078),
            .ce(),
            .sr(N__48625));
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_8_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_8_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__27271),
            .in2(N__27275),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_8_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_8_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(N__26930),
            .in2(N__26918),
            .in3(N__25064),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_8_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_8_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(N__27281),
            .in2(N__27065),
            .in3(N__25061),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_8_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_8_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(N__27227),
            .in2(N__27290),
            .in3(N__25058),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_8_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_8_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__25055),
            .in2(N__25046),
            .in3(N__25022),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(N__25202),
            .in2(N__27167),
            .in3(N__25187),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(N__25184),
            .in2(N__27113),
            .in3(N__25160),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_16_7  (
            .in0(_gnd_net_),
            .in1(N__27959),
            .in2(N__27887),
            .in3(N__25157),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__25154),
            .in2(N__25148),
            .in3(N__25130),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__25127),
            .in2(N__27476),
            .in3(N__25109),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__27644),
            .in2(N__27221),
            .in3(N__25106),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__28070),
            .in2(N__27452),
            .in3(N__25103),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__41225),
            .in2(N__27443),
            .in3(N__25091),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__25088),
            .in2(N__27380),
            .in3(N__25067),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__27467),
            .in2(N__29867),
            .in3(N__25340),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__27767),
            .in2(N__27461),
            .in3(N__25328),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__25325),
            .in2(N__27653),
            .in3(N__25304),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__29777),
            .in2(N__27584),
            .in3(N__25292),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__25289),
            .in2(N__27323),
            .in3(N__25268),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__25265),
            .in2(N__27593),
            .in3(N__25241),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__35420),
            .in2(N__27308),
            .in3(N__25226),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__25223),
            .in2(N__27704),
            .in3(N__25205),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__27536),
            .in2(N__27761),
            .in3(N__25427),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__29945),
            .in2(N__27899),
            .in3(N__25418),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__29852),
            .in2(N__29708),
            .in3(N__25406),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__25523),
            .in2(N__28022),
            .in3(N__25403),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__25511),
            .in2(N__27968),
            .in3(N__25391),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__25517),
            .in2(N__27908),
            .in3(N__25379),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__25376),
            .in2(N__30041),
            .in3(N__25361),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__25460),
            .in2(N__30316),
            .in3(N__25352),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__30312),
            .in2(N__42710),
            .in3(N__25541),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__25538),
            .in2(N__30317),
            .in3(N__25529),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_0  (
            .in0(N__35402),
            .in1(N__31922),
            .in2(_gnd_net_),
            .in3(N__25526),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_8_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_8_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28043),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27931),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27994),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_8_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_8_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25487),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_8_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_8_21_1 .LUT_INIT=16'b0010001011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_8_21_1  (
            .in0(N__31992),
            .in1(N__32397),
            .in2(N__32224),
            .in3(N__25454),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49036),
            .ce(),
            .sr(N__48655));
    defparam \phase_controller_inst2.S2_LC_8_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_8_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_8_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26996),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49036),
            .ce(),
            .sr(N__48655));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_9_4_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_9_4_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_9_4_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_9_4_0  (
            .in0(N__25942),
            .in1(N__25776),
            .in2(_gnd_net_),
            .in3(N__25568),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__49143),
            .ce(N__25829),
            .sr(N__48527));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_9_4_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_9_4_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_9_4_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_9_4_1  (
            .in0(N__25938),
            .in1(N__25749),
            .in2(_gnd_net_),
            .in3(N__25565),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__49143),
            .ce(N__25829),
            .sr(N__48527));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_9_4_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_9_4_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_9_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_9_4_2  (
            .in0(N__25943),
            .in1(N__25726),
            .in2(_gnd_net_),
            .in3(N__25562),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__49143),
            .ce(N__25829),
            .sr(N__48527));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_9_4_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_9_4_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_9_4_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_9_4_3  (
            .in0(N__25939),
            .in1(N__25698),
            .in2(_gnd_net_),
            .in3(N__25559),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__49143),
            .ce(N__25829),
            .sr(N__48527));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_9_4_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_9_4_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_9_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_9_4_4  (
            .in0(N__25944),
            .in1(N__25668),
            .in2(_gnd_net_),
            .in3(N__25556),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__49143),
            .ce(N__25829),
            .sr(N__48527));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_9_4_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_9_4_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_9_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_9_4_5  (
            .in0(N__25940),
            .in1(N__25641),
            .in2(_gnd_net_),
            .in3(N__25553),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__49143),
            .ce(N__25829),
            .sr(N__48527));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_9_4_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_9_4_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_9_4_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_9_4_6  (
            .in0(N__25945),
            .in1(N__26161),
            .in2(_gnd_net_),
            .in3(N__25550),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__49143),
            .ce(N__25829),
            .sr(N__48527));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_9_4_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_9_4_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_9_4_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_9_4_7  (
            .in0(N__25941),
            .in1(N__26137),
            .in2(_gnd_net_),
            .in3(N__25547),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__49143),
            .ce(N__25829),
            .sr(N__48527));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_9_5_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_9_5_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_9_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_9_5_0  (
            .in0(N__25927),
            .in1(N__26106),
            .in2(_gnd_net_),
            .in3(N__25544),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__49139),
            .ce(N__25818),
            .sr(N__48531));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_9_5_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_9_5_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_9_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_9_5_1  (
            .in0(N__25931),
            .in1(N__26079),
            .in2(_gnd_net_),
            .in3(N__25595),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__49139),
            .ce(N__25818),
            .sr(N__48531));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_9_5_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_9_5_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_9_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_9_5_2  (
            .in0(N__25924),
            .in1(N__26050),
            .in2(_gnd_net_),
            .in3(N__25592),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__49139),
            .ce(N__25818),
            .sr(N__48531));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_9_5_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_9_5_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_9_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_9_5_3  (
            .in0(N__25928),
            .in1(N__26022),
            .in2(_gnd_net_),
            .in3(N__25589),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__49139),
            .ce(N__25818),
            .sr(N__48531));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_9_5_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_9_5_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_9_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_9_5_4  (
            .in0(N__25925),
            .in1(N__25995),
            .in2(_gnd_net_),
            .in3(N__25586),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__49139),
            .ce(N__25818),
            .sr(N__48531));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_9_5_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_9_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_9_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_9_5_5  (
            .in0(N__25929),
            .in1(N__25974),
            .in2(_gnd_net_),
            .in3(N__25583),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__49139),
            .ce(N__25818),
            .sr(N__48531));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_9_5_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_9_5_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_9_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_9_5_6  (
            .in0(N__25926),
            .in1(N__26392),
            .in2(_gnd_net_),
            .in3(N__25580),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__49139),
            .ce(N__25818),
            .sr(N__48531));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_9_5_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_9_5_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_9_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_9_5_7  (
            .in0(N__25930),
            .in1(N__26367),
            .in2(_gnd_net_),
            .in3(N__25577),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__49139),
            .ce(N__25818),
            .sr(N__48531));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_9_6_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_9_6_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_9_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_9_6_0  (
            .in0(N__25920),
            .in1(N__26334),
            .in2(_gnd_net_),
            .in3(N__25574),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__49136),
            .ce(N__25809),
            .sr(N__48538));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_9_6_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_9_6_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_9_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_9_6_1  (
            .in0(N__25946),
            .in1(N__26307),
            .in2(_gnd_net_),
            .in3(N__25571),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__49136),
            .ce(N__25809),
            .sr(N__48538));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_9_6_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_9_6_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_9_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_9_6_2  (
            .in0(N__25921),
            .in1(N__26283),
            .in2(_gnd_net_),
            .in3(N__25622),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__49136),
            .ce(N__25809),
            .sr(N__48538));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_9_6_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_9_6_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_9_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_9_6_3  (
            .in0(N__25947),
            .in1(N__26262),
            .in2(_gnd_net_),
            .in3(N__25619),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__49136),
            .ce(N__25809),
            .sr(N__48538));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_9_6_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_9_6_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_9_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_9_6_4  (
            .in0(N__25922),
            .in1(N__26235),
            .in2(_gnd_net_),
            .in3(N__25616),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__49136),
            .ce(N__25809),
            .sr(N__48538));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_9_6_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_9_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_9_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_9_6_5  (
            .in0(N__25948),
            .in1(N__26208),
            .in2(_gnd_net_),
            .in3(N__25613),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__49136),
            .ce(N__25809),
            .sr(N__48538));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_9_6_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_9_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_9_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_9_6_6  (
            .in0(N__25923),
            .in1(N__26182),
            .in2(_gnd_net_),
            .in3(N__25610),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__49136),
            .ce(N__25809),
            .sr(N__48538));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_9_6_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_9_6_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_9_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_9_6_7  (
            .in0(N__25949),
            .in1(N__26658),
            .in2(_gnd_net_),
            .in3(N__25607),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__49136),
            .ce(N__25809),
            .sr(N__48538));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_9_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_9_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_9_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_9_7_0  (
            .in0(N__25932),
            .in1(N__26625),
            .in2(_gnd_net_),
            .in3(N__25604),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__49132),
            .ce(N__25825),
            .sr(N__48544));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_9_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_9_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_9_7_1  (
            .in0(N__25936),
            .in1(N__26601),
            .in2(_gnd_net_),
            .in3(N__25601),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__49132),
            .ce(N__25825),
            .sr(N__48544));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_9_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_9_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_9_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_9_7_2  (
            .in0(N__25933),
            .in1(N__26577),
            .in2(_gnd_net_),
            .in3(N__25598),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__49132),
            .ce(N__25825),
            .sr(N__48544));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_9_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_9_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_9_7_3  (
            .in0(N__25937),
            .in1(N__26517),
            .in2(_gnd_net_),
            .in3(N__25955),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__49132),
            .ce(N__25825),
            .sr(N__48544));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_9_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_9_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_9_7_4  (
            .in0(N__25934),
            .in1(N__26557),
            .in2(_gnd_net_),
            .in3(N__25952),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__49132),
            .ce(N__25825),
            .sr(N__48544));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_9_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_9_7_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_9_7_5  (
            .in0(N__26536),
            .in1(N__25935),
            .in2(_gnd_net_),
            .in3(N__25832),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49132),
            .ce(N__25825),
            .sr(N__48544));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_8_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__25732),
            .in2(N__25787),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49127),
            .ce(N__26490),
            .sr(N__48551));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__25756),
            .in2(N__25709),
            .in3(N__25736),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49127),
            .ce(N__26490),
            .sr(N__48551));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__25733),
            .in2(N__25675),
            .in3(N__25712),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49127),
            .ce(N__26490),
            .sr(N__48551));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__25708),
            .in2(N__25648),
            .in3(N__25679),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49127),
            .ce(N__26490),
            .sr(N__48551));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__26167),
            .in2(N__25676),
            .in3(N__25652),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49127),
            .ce(N__26490),
            .sr(N__48551));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__26143),
            .in2(N__25649),
            .in3(N__25625),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49127),
            .ce(N__26490),
            .sr(N__48551));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__26168),
            .in2(N__26119),
            .in3(N__26147),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49127),
            .ce(N__26490),
            .sr(N__48551));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__26144),
            .in2(N__26086),
            .in3(N__26123),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49127),
            .ce(N__26490),
            .sr(N__48551));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__26056),
            .in2(N__26120),
            .in3(N__26090),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49121),
            .ce(N__26483),
            .sr(N__48559));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__26029),
            .in2(N__26087),
            .in3(N__26060),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49121),
            .ce(N__26483),
            .sr(N__48559));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__26057),
            .in2(N__26002),
            .in3(N__26036),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49121),
            .ce(N__26483),
            .sr(N__48559));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__25975),
            .in2(N__26033),
            .in3(N__26006),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49121),
            .ce(N__26483),
            .sr(N__48559));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__26398),
            .in2(N__26003),
            .in3(N__25979),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49121),
            .ce(N__26483),
            .sr(N__48559));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__25976),
            .in2(N__26374),
            .in3(N__25958),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49121),
            .ce(N__26483),
            .sr(N__48559));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__26399),
            .in2(N__26347),
            .in3(N__26378),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49121),
            .ce(N__26483),
            .sr(N__48559));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__26308),
            .in2(N__26375),
            .in3(N__26351),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49121),
            .ce(N__26483),
            .sr(N__48559));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__26284),
            .in2(N__26348),
            .in3(N__26318),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49113),
            .ce(N__26491),
            .sr(N__48572));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__26263),
            .in2(N__26315),
            .in3(N__26288),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49113),
            .ce(N__26491),
            .sr(N__48572));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__26285),
            .in2(N__26242),
            .in3(N__26267),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49113),
            .ce(N__26491),
            .sr(N__48572));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__26264),
            .in2(N__26215),
            .in3(N__26246),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49113),
            .ce(N__26491),
            .sr(N__48572));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__26188),
            .in2(N__26243),
            .in3(N__26219),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49113),
            .ce(N__26491),
            .sr(N__48572));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__26665),
            .in2(N__26216),
            .in3(N__26192),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49113),
            .ce(N__26491),
            .sr(N__48572));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__26189),
            .in2(N__26638),
            .in3(N__26672),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49113),
            .ce(N__26491),
            .sr(N__48572));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__26602),
            .in2(N__26669),
            .in3(N__26642),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49113),
            .ce(N__26491),
            .sr(N__48572));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__26578),
            .in2(N__26639),
            .in3(N__26609),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49105),
            .ce(N__26492),
            .sr(N__48582));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__26518),
            .in2(N__26606),
            .in3(N__26582),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49105),
            .ce(N__26492),
            .sr(N__48582));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__26579),
            .in2(N__26561),
            .in3(N__26543),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49105),
            .ce(N__26492),
            .sr(N__48582));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__26540),
            .in2(N__26522),
            .in3(N__26498),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49105),
            .ce(N__26492),
            .sr(N__48582));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26495),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49105),
            .ce(N__26492),
            .sr(N__48582));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_12_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_12_0  (
            .in0(N__26423),
            .in1(N__26443),
            .in2(_gnd_net_),
            .in3(N__34701),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_9_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_9_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_9_12_1 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_27_LC_9_12_1  (
            .in0(N__34702),
            .in1(N__26424),
            .in2(N__26402),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49097),
            .ce(N__34242),
            .sr(N__48589));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_12_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_12_2  (
            .in0(N__26864),
            .in1(N__26890),
            .in2(_gnd_net_),
            .in3(N__34700),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_9_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_9_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_9_12_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_28_LC_9_12_3  (
            .in0(N__34703),
            .in1(_gnd_net_),
            .in2(N__26879),
            .in3(N__26865),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49097),
            .ce(N__34242),
            .sr(N__48589));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_4 .LUT_INIT=16'b1011001010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_4  (
            .in0(N__26803),
            .in1(N__30931),
            .in2(N__26843),
            .in3(N__30538),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_12_5 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_12_5  (
            .in0(N__30932),
            .in1(N__26804),
            .in2(N__30539),
            .in3(N__26842),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_9_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_9_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_9_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_29_LC_9_12_6  (
            .in0(N__26831),
            .in1(N__28547),
            .in2(_gnd_net_),
            .in3(N__34704),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49097),
            .ce(N__34242),
            .sr(N__48589));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_12_7 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_12_7  (
            .in0(N__29405),
            .in1(N__30563),
            .in2(N__30596),
            .in3(N__29393),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_9_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_9_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_9_13_0 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst2.state_0_LC_9_13_0  (
            .in0(N__26988),
            .in1(N__27033),
            .in2(N__26693),
            .in3(N__26705),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49088),
            .ce(),
            .sr(N__48600));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_9_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_9_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_9_13_1 .LUT_INIT=16'b1000110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_9_13_1  (
            .in0(N__26704),
            .in1(N__26791),
            .in2(N__26765),
            .in3(N__26736),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49088),
            .ce(),
            .sr(N__48600));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_9_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_9_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__26703),
            .in2(_gnd_net_),
            .in3(N__26689),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(\phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_3_LC_9_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_9_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_9_13_3 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst2.state_3_LC_9_13_3  (
            .in0(N__31649),
            .in1(N__31681),
            .in2(N__27056),
            .in3(N__33659),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49088),
            .ce(),
            .sr(N__48600));
    defparam \phase_controller_inst2.state_2_LC_9_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_9_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_9_13_5 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst2.state_2_LC_9_13_5  (
            .in0(N__27049),
            .in1(N__31680),
            .in2(N__35744),
            .in3(N__31650),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49088),
            .ce(),
            .sr(N__48600));
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_9_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_9_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNIG7JF_2_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__27048),
            .in2(_gnd_net_),
            .in3(N__35739),
            .lcout(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ),
            .ltout(\phase_controller_inst2.state_RNIG7JFZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_1_LC_9_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_9_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_9_13_7 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \phase_controller_inst2.state_1_LC_9_13_7  (
            .in0(N__27034),
            .in1(_gnd_net_),
            .in2(N__26999),
            .in3(N__26989),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49088),
            .ce(),
            .sr(N__48600));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_14_0 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_9_14_0  (
            .in0(N__32390),
            .in1(N__32154),
            .in2(_gnd_net_),
            .in3(N__26969),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49079),
            .ce(),
            .sr(N__48608));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_9_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_9_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33006),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26941),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_0 ),
            .ltout(\current_shift_inst.PI_CTRL.integrator_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_9_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_9_14_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_9_14_3  (
            .in0(N__35292),
            .in1(N__33007),
            .in2(N__26921),
            .in3(N__29351),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_14_4 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_9_14_4  (
            .in0(N__32391),
            .in1(N__32155),
            .in2(_gnd_net_),
            .in3(N__26903),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49079),
            .ce(),
            .sr(N__48608));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_14_7 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_9_14_7  (
            .in0(N__32153),
            .in1(N__32392),
            .in2(_gnd_net_),
            .in3(N__27299),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49079),
            .ce(),
            .sr(N__48608));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_9_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_9_15_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_9_15_0  (
            .in0(N__35336),
            .in1(N__27241),
            .in2(N__33886),
            .in3(N__29543),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27083),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_9_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_9_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_9_15_2  (
            .in0(N__35334),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_9_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_9_15_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_9_15_3  (
            .in0(N__27240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_9_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_9_15_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_9_15_4  (
            .in0(N__35339),
            .in1(N__31857),
            .in2(N__33299),
            .in3(N__29456),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_9_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_9_15_5 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_9_15_5  (
            .in0(N__27201),
            .in1(N__35337),
            .in2(N__29522),
            .in3(N__33964),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_9_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_9_15_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_9_15_6  (
            .in0(N__35338),
            .in1(N__27157),
            .in2(N__33482),
            .in3(N__29510),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_9_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_9_15_7 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_9_15_7  (
            .in0(N__33923),
            .in1(N__35335),
            .in2(N__29342),
            .in3(N__27084),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_9_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_9_16_0 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_9_16_0  (
            .in0(N__33188),
            .in1(N__27528),
            .in2(N__35397),
            .in3(N__29465),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_9_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_9_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33187),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_9_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_9_16_2 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_9_16_2  (
            .in0(N__29909),
            .in1(N__35354),
            .in2(N__33416),
            .in3(N__29603),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_9_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_9_16_3 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_9_16_3  (
            .in0(N__27818),
            .in1(N__35368),
            .in2(N__31469),
            .in3(N__29594),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_9_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_9_16_4 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_9_16_4  (
            .in0(N__28234),
            .in1(N__29630),
            .in2(N__35398),
            .in3(N__33347),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_9_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_9_16_5 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_9_16_5  (
            .in0(N__41276),
            .in1(N__33323),
            .in2(N__35395),
            .in3(N__29621),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_9_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_9_16_6 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_9_16_6  (
            .in0(N__27409),
            .in1(N__33440),
            .in2(N__35399),
            .in3(N__29612),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_9_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_9_16_7 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_9_16_7  (
            .in0(N__27352),
            .in1(N__35129),
            .in2(N__35396),
            .in3(N__29561),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_9_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_9_17_0 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_9_17_0  (
            .in0(N__35461),
            .in1(N__30024),
            .in2(N__35384),
            .in3(N__29696),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27808),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_9_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_9_17_2 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_9_17_2  (
            .in0(N__27575),
            .in1(N__31418),
            .in2(N__35383),
            .in3(N__29678),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_9_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_9_17_3 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_9_17_3  (
            .in0(N__27748),
            .in1(N__35330),
            .in2(N__32435),
            .in3(N__29687),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_9_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_9_17_4 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_9_17_4  (
            .in0(N__27694),
            .in1(N__32459),
            .in2(N__35381),
            .in3(N__29585),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_9_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_9_17_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_9_17_5  (
            .in0(N__31843),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_9_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_9_17_6 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_9_17_6  (
            .in0(N__27634),
            .in1(N__32483),
            .in2(N__35382),
            .in3(N__29552),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_9_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_9_17_7 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_9_17_7  (
            .in0(N__31493),
            .in1(N__29839),
            .in2(N__29576),
            .in3(N__35320),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_9_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_9_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27567),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28205),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_9_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_9_18_3 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_9_18_3  (
            .in0(N__31445),
            .in1(N__28052),
            .in2(N__35401),
            .in3(N__29657),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_9_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_9_18_4 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_9_18_4  (
            .in0(N__28013),
            .in1(N__35375),
            .in2(N__29936),
            .in3(N__29648),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_18_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_18_5  (
            .in0(N__27837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_9_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_9_18_6 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_9_18_6  (
            .in0(N__27949),
            .in1(N__35376),
            .in2(N__30005),
            .in3(N__29639),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_9_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_9_18_7 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_9_18_7  (
            .in0(N__32507),
            .in1(N__29977),
            .in2(N__35400),
            .in3(N__29669),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_9_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_9_19_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_9_19_0  (
            .in0(N__27854),
            .in1(N__33389),
            .in2(N__35403),
            .in3(N__29501),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_9_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_9_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_9_19_2 .LUT_INIT=16'b0000000111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_9_19_2  (
            .in0(N__31947),
            .in1(N__32389),
            .in2(N__32215),
            .in3(N__27875),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49046),
            .ce(),
            .sr(N__48641));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_9_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_9_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_9_19_4 .LUT_INIT=16'b0010001011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_9_19_4  (
            .in0(N__31945),
            .in1(N__32387),
            .in2(N__32213),
            .in3(N__27824),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49046),
            .ce(),
            .sr(N__48641));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_9_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_9_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_9_19_5 .LUT_INIT=16'b0100111101001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_9_19_5  (
            .in0(N__32386),
            .in1(N__31949),
            .in2(N__28319),
            .in3(N__32188),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49046),
            .ce(),
            .sr(N__48641));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_9_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_9_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_9_19_6 .LUT_INIT=16'b0010001011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_9_19_6  (
            .in0(N__31946),
            .in1(N__32388),
            .in2(N__32214),
            .in3(N__28307),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49046),
            .ce(),
            .sr(N__48641));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_9_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_9_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_9_19_7 .LUT_INIT=16'b0100111101001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_9_19_7  (
            .in0(N__32385),
            .in1(N__31948),
            .in2(N__28253),
            .in3(N__32187),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49046),
            .ce(),
            .sr(N__48641));
    defparam \delay_measurement_inst.stop_timer_tr_LC_9_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_9_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_9_20_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_9_20_0  (
            .in0(N__28135),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28118),
            .ce(),
            .sr(N__48646));
    defparam \delay_measurement_inst.start_timer_tr_LC_9_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_9_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_9_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28134),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28118),
            .ce(),
            .sr(N__48646));
    defparam \phase_controller_inst2.S1_LC_9_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31654),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49017),
            .ce(),
            .sr(N__48658));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6 (
            .in0(N__28100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_10_4_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_10_4_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_10_4_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_10_4_4 (
            .in0(N__28082),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49137),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_5_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_5_4  (
            .in0(N__30238),
            .in1(N__30273),
            .in2(_gnd_net_),
            .in3(N__34532),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_10_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_10_7_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__30368),
            .in2(_gnd_net_),
            .in3(N__30113),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_10_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_10_7_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_10_7_2  (
            .in0(N__28454),
            .in1(N__30263),
            .in2(N__28478),
            .in3(N__28361),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_7_3 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_7_3  (
            .in0(N__28475),
            .in1(N__28748),
            .in2(N__28466),
            .in3(N__28520),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_4  (
            .in0(N__28455),
            .in1(_gnd_net_),
            .in2(N__28436),
            .in3(N__28429),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49122),
            .ce(N__34199),
            .sr(N__48532));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0  (
            .in0(N__34468),
            .in1(N__28381),
            .in2(_gnd_net_),
            .in3(N__28399),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__28380),
            .in2(N__28388),
            .in3(N__34472),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49114),
            .ce(N__34183),
            .sr(N__48539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_8_4  (
            .in0(N__28379),
            .in1(N__32630),
            .in2(N__28605),
            .in3(N__28334),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5  (
            .in0(N__28335),
            .in1(N__28351),
            .in2(_gnd_net_),
            .in3(N__34469),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(elapsed_time_ns_1_RNILK91B_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6  (
            .in0(N__34470),
            .in1(_gnd_net_),
            .in2(N__28340),
            .in3(N__28336),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49114),
            .ce(N__34183),
            .sr(N__48539));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_10_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_10_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_10_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_10_8_7  (
            .in0(N__28604),
            .in1(N__34471),
            .in2(_gnd_net_),
            .in3(N__28580),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49114),
            .ce(N__34183),
            .sr(N__48539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_10_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_10_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_10_9_0  (
            .in0(N__28793),
            .in1(N__29433),
            .in2(N__28557),
            .in3(N__29124),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_10_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_10_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_10_9_1  (
            .in0(N__28499),
            .in1(N__28505),
            .in2(N__28523),
            .in3(N__28511),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_10_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_10_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_10_9_2  (
            .in0(N__28649),
            .in1(N__32838),
            .in2(N__32805),
            .in3(N__28673),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_10_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_10_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_10_9_3  (
            .in0(N__29003),
            .in1(N__28938),
            .in2(N__32922),
            .in3(N__28884),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_10_9_4  (
            .in0(N__30180),
            .in1(N__29067),
            .in2(N__32700),
            .in3(N__34724),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_7  (
            .in0(N__28629),
            .in1(N__28650),
            .in2(_gnd_net_),
            .in3(N__34598),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_10_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_10_10_0 .LUT_INIT=16'b0010101100001010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_10_10_0  (
            .in0(N__30880),
            .in1(N__30906),
            .in2(N__28720),
            .in3(N__28702),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_10_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_10_1  (
            .in0(N__28790),
            .in1(N__34511),
            .in2(_gnd_net_),
            .in3(N__28489),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_2  (
            .in0(N__34513),
            .in1(_gnd_net_),
            .in2(N__28796),
            .in3(N__28791),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49098),
            .ce(N__34259),
            .sr(N__48552));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_10_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_10_3  (
            .in0(N__28742),
            .in1(_gnd_net_),
            .in2(N__28768),
            .in3(N__34512),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(elapsed_time_ns_1_RNI0CQBB_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_10_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_10_10_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_31_LC_10_10_4  (
            .in0(N__34514),
            .in1(_gnd_net_),
            .in2(N__28751),
            .in3(N__28743),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49098),
            .ce(N__34259),
            .sr(N__48552));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_10_5 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_10_5  (
            .in0(N__28703),
            .in1(N__28719),
            .in2(N__30911),
            .in3(N__30881),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_10_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_10_10_6 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_10_10_6  (
            .in0(N__30879),
            .in1(N__30907),
            .in2(N__28721),
            .in3(N__28701),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_10_10_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_10_10_7  (
            .in0(N__28691),
            .in1(N__34515),
            .in2(_gnd_net_),
            .in3(N__28676),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49098),
            .ce(N__34259),
            .sr(N__48552));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0  (
            .in0(N__30475),
            .in1(N__30492),
            .in2(N__28985),
            .in3(N__28925),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_10_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_10_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_10_11_2  (
            .in0(N__28655),
            .in1(N__28630),
            .in2(_gnd_net_),
            .in3(N__34591),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49090),
            .ce(N__34250),
            .sr(N__48563));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_3 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_3  (
            .in0(N__28924),
            .in1(N__30474),
            .in2(N__30497),
            .in3(N__28981),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_11_4  (
            .in0(N__29004),
            .in1(N__29026),
            .in2(_gnd_net_),
            .in3(N__34588),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_10_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_10_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_10_11_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_10_11_5  (
            .in0(N__34590),
            .in1(_gnd_net_),
            .in2(N__29015),
            .in3(N__29005),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49090),
            .ce(N__34250),
            .sr(N__48563));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_11_6  (
            .in0(N__28947),
            .in1(N__28966),
            .in2(_gnd_net_),
            .in3(N__34587),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_10_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_10_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_10_11_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_10_11_7  (
            .in0(N__34589),
            .in1(_gnd_net_),
            .in2(N__28955),
            .in3(N__28948),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49090),
            .ce(N__34250),
            .sr(N__48563));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_12_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_12_0  (
            .in0(N__30456),
            .in1(N__28868),
            .in2(N__34274),
            .in3(N__30702),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_1  (
            .in0(N__28893),
            .in1(N__28909),
            .in2(_gnd_net_),
            .in3(N__34592),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_10_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_10_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_10_12_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_20_LC_10_12_2  (
            .in0(N__34594),
            .in1(_gnd_net_),
            .in2(N__28898),
            .in3(N__28894),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49081),
            .ce(N__34244),
            .sr(N__48573));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_12_3 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_12_3  (
            .in0(N__28867),
            .in1(N__34273),
            .in2(N__30707),
            .in3(N__30457),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_10_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_10_12_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_10_12_4  (
            .in0(N__34593),
            .in1(N__28859),
            .in2(_gnd_net_),
            .in3(N__28829),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49081),
            .ce(N__34244),
            .sr(N__48573));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_10_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_10_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_10_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_10_12_5  (
            .in0(N__29330),
            .in1(N__29303),
            .in2(_gnd_net_),
            .in3(N__34596),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49081),
            .ce(N__34244),
            .sr(N__48573));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_10_12_6  (
            .in0(N__34595),
            .in1(N__29270),
            .in2(_gnd_net_),
            .in3(N__29243),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49081),
            .ce(N__34244),
            .sr(N__48573));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_10_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_10_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_10_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_10_12_7  (
            .in0(N__29216),
            .in1(N__29189),
            .in2(_gnd_net_),
            .in3(N__34597),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49081),
            .ce(N__34244),
            .sr(N__48573));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_13_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_13_0  (
            .in0(N__29044),
            .in1(N__30615),
            .in2(N__29105),
            .in3(N__30638),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_13_1 .LUT_INIT=16'b1111011100110001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_13_1  (
            .in0(N__30637),
            .in1(N__30616),
            .in2(N__29048),
            .in3(N__29101),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_13_2  (
            .in0(N__34602),
            .in1(N__29139),
            .in2(_gnd_net_),
            .in3(N__29152),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_10_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_10_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_10_13_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_25_LC_10_13_3  (
            .in0(N__29140),
            .in1(_gnd_net_),
            .in2(N__29108),
            .in3(N__34605),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49071),
            .ce(N__34245),
            .sr(N__48583));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_13_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_13_4  (
            .in0(N__29074),
            .in1(_gnd_net_),
            .in2(N__34684),
            .in3(N__29086),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(elapsed_time_ns_1_RNI2DPBB_0_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_10_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_10_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_10_13_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_24_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__29075),
            .in2(N__29051),
            .in3(N__34604),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49071),
            .ce(N__34245),
            .sr(N__48583));
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_10_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_10_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_10_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_26_LC_10_13_6  (
            .in0(N__34603),
            .in1(N__29445),
            .in2(_gnd_net_),
            .in3(N__29420),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49071),
            .ce(N__34245),
            .sr(N__48583));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_13_7 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_13_7  (
            .in0(N__29404),
            .in1(N__30558),
            .in2(N__30592),
            .in3(N__29392),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_10_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_10_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__29381),
            .in2(_gnd_net_),
            .in3(N__33715),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_10_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_10_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__29375),
            .in2(_gnd_net_),
            .in3(N__33088),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_10_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_10_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__29369),
            .in2(_gnd_net_),
            .in3(N__33052),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_10_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_10_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__29363),
            .in2(_gnd_net_),
            .in3(N__33155),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_10_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_10_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__29357),
            .in2(_gnd_net_),
            .in3(N__29345),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_10_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_10_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__33896),
            .in2(_gnd_net_),
            .in3(N__29333),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_10_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_10_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__33851),
            .in2(_gnd_net_),
            .in3(N__29537),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_10_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_10_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__33812),
            .in2(_gnd_net_),
            .in3(N__29525),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_10_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_10_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__33935),
            .in2(_gnd_net_),
            .in3(N__29513),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_8 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_10_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_10_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__33449),
            .in2(_gnd_net_),
            .in3(N__29504),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_10_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_10_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__33356),
            .in2(_gnd_net_),
            .in3(N__29489),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_10_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_10_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__33491),
            .in2(_gnd_net_),
            .in3(N__29474),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_10_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_10_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__29471),
            .in2(_gnd_net_),
            .in3(N__29459),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_10_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_10_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__33266),
            .in2(_gnd_net_),
            .in3(N__29450),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_10_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_10_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__33343),
            .in2(_gnd_net_),
            .in3(N__29624),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_10_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_10_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__33319),
            .in2(_gnd_net_),
            .in3(N__29615),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_10_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_10_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__33439),
            .in2(_gnd_net_),
            .in3(N__29606),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_10_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_10_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__33412),
            .in2(_gnd_net_),
            .in3(N__29597),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_10_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_10_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__31461),
            .in2(_gnd_net_),
            .in3(N__29588),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_10_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_10_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__32451),
            .in2(_gnd_net_),
            .in3(N__29579),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_10_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_10_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__31485),
            .in2(_gnd_net_),
            .in3(N__29564),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_10_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_10_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__35128),
            .in2(_gnd_net_),
            .in3(N__29555),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_10_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_10_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__32475),
            .in2(_gnd_net_),
            .in3(N__29546),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_10_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_10_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__30026),
            .in2(_gnd_net_),
            .in3(N__29690),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_10_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_10_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__32424),
            .in2(_gnd_net_),
            .in3(N__29681),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_10_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_10_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__31410),
            .in2(_gnd_net_),
            .in3(N__29672),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_10_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_10_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__32499),
            .in2(_gnd_net_),
            .in3(N__29663),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_10_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_10_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__33637),
            .in2(_gnd_net_),
            .in3(N__29660),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_10_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_10_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31441),
            .in3(N__29651),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_10_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_10_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__29931),
            .in2(_gnd_net_),
            .in3(N__29642),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_10_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_10_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__30000),
            .in2(_gnd_net_),
            .in3(N__29633),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_10_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_10_17_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_10_17_7  (
            .in0(N__30094),
            .in1(N__35358),
            .in2(_gnd_net_),
            .in3(N__30044),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__30025),
            .in2(_gnd_net_),
            .in3(N__35331),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_18_2  (
            .in0(N__30004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35333),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_10_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_10_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29976),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_10_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_10_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_10_18_4  (
            .in0(N__29935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35332),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_10_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_10_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29908),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29755),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_10_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_10_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29824),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_10_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_10_19_2 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_10_19_2  (
            .in0(N__33641),
            .in1(N__29768),
            .in2(N__35404),
            .in3(N__29717),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_10_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_10_19_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_10_19_4  (
            .in0(N__35391),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_11_4_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_11_4_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_11_4_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_11_4_3 (
            .in0(N__30296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49133),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_11_4_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_11_4_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_11_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_11_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30284),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49133),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_11_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_11_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_11_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_11_5_7  (
            .in0(N__30278),
            .in1(N__30234),
            .in2(_gnd_net_),
            .in3(N__34606),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49129),
            .ce(N__34251),
            .sr(N__48521));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0  (
            .in0(N__30659),
            .in1(N__30682),
            .in2(N__30164),
            .in3(N__32672),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_1  (
            .in0(N__32671),
            .in1(N__30658),
            .in2(N__30686),
            .in3(N__30160),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_7_2  (
            .in0(N__30195),
            .in1(N__34575),
            .in2(_gnd_net_),
            .in3(N__30211),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(elapsed_time_ns_1_RNI1CPBB_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_11_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_11_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_11_7_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_23_LC_11_7_3  (
            .in0(N__34576),
            .in1(_gnd_net_),
            .in2(N__30200),
            .in3(N__30196),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49115),
            .ce(N__34243),
            .sr(N__48528));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_11_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_11_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_11_7_6  (
            .in0(N__30152),
            .in1(N__30131),
            .in2(_gnd_net_),
            .in3(N__34578),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49115),
            .ce(N__34243),
            .sr(N__48528));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_11_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_11_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_11_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_11_7_7  (
            .in0(N__34577),
            .in1(N__30404),
            .in2(_gnd_net_),
            .in3(N__30383),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49115),
            .ce(N__34243),
            .sr(N__48528));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_11_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_11_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_11_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35099),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49107),
            .ce(),
            .sr(N__48533));
    defparam \phase_controller_inst1.stoper_tr.running_LC_11_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_11_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_11_8_3 .LUT_INIT=16'b1011101000111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_11_8_3  (
            .in0(N__30338),
            .in1(N__34962),
            .in2(N__34941),
            .in3(N__35003),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49107),
            .ce(),
            .sr(N__48533));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_11_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_11_8_4 .LUT_INIT=16'b1111110101110101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_11_8_4  (
            .in0(N__34961),
            .in1(N__30350),
            .in2(N__31531),
            .in3(N__31511),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_11_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_11_8_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30341),
            .in3(N__34925),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_8_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_8_6  (
            .in0(N__34960),
            .in1(N__30337),
            .in2(_gnd_net_),
            .in3(N__35098),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_11_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_11_8_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30329),
            .in3(N__30856),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__30326),
            .in2(N__30839),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_9_1  (
            .in0(N__34175),
            .in1(N__30793),
            .in2(_gnd_net_),
            .in3(N__30320),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49099),
            .ce(),
            .sr(N__48540));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_9_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_9_2  (
            .in0(N__34252),
            .in1(N__30766),
            .in2(N__30440),
            .in3(N__30431),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49099),
            .ce(),
            .sr(N__48540));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_9_3  (
            .in0(N__34176),
            .in1(N__30727),
            .in2(_gnd_net_),
            .in3(N__30428),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49099),
            .ce(),
            .sr(N__48540));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_9_4  (
            .in0(N__34253),
            .in1(N__31186),
            .in2(_gnd_net_),
            .in3(N__30425),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49099),
            .ce(),
            .sr(N__48540));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_9_5  (
            .in0(N__34177),
            .in1(N__31147),
            .in2(_gnd_net_),
            .in3(N__30422),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49099),
            .ce(),
            .sr(N__48540));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_9_6  (
            .in0(N__34254),
            .in1(N__31096),
            .in2(_gnd_net_),
            .in3(N__30419),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49099),
            .ce(),
            .sr(N__48540));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_9_7  (
            .in0(N__34178),
            .in1(N__31057),
            .in2(_gnd_net_),
            .in3(N__30416),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49099),
            .ce(),
            .sr(N__48540));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_10_0  (
            .in0(N__34182),
            .in1(N__31018),
            .in2(_gnd_net_),
            .in3(N__30413),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49091),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_10_1  (
            .in0(N__34163),
            .in1(N__30994),
            .in2(_gnd_net_),
            .in3(N__30410),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49091),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_10_2  (
            .in0(N__34179),
            .in1(N__30955),
            .in2(_gnd_net_),
            .in3(N__30407),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49091),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_10_3  (
            .in0(N__34164),
            .in1(N__31378),
            .in2(_gnd_net_),
            .in3(N__30515),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49091),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_10_4  (
            .in0(N__34180),
            .in1(N__31357),
            .in2(_gnd_net_),
            .in3(N__30512),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49091),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_10_5  (
            .in0(N__34165),
            .in1(N__31318),
            .in2(_gnd_net_),
            .in3(N__30509),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49091),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_10_6  (
            .in0(N__34181),
            .in1(N__31294),
            .in2(_gnd_net_),
            .in3(N__30506),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49091),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_10_7  (
            .in0(N__34166),
            .in1(N__32564),
            .in2(_gnd_net_),
            .in3(N__30503),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49091),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_11_0  (
            .in0(N__34246),
            .in1(N__32584),
            .in2(_gnd_net_),
            .in3(N__30500),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49082),
            .ce(),
            .sr(N__48553));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_11_1  (
            .in0(N__34189),
            .in1(N__30496),
            .in2(_gnd_net_),
            .in3(N__30479),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49082),
            .ce(),
            .sr(N__48553));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_11_2  (
            .in0(N__34247),
            .in1(N__30476),
            .in2(_gnd_net_),
            .in3(N__30461),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49082),
            .ce(),
            .sr(N__48553));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_11_3  (
            .in0(N__34190),
            .in1(N__30458),
            .in2(_gnd_net_),
            .in3(N__30443),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49082),
            .ce(),
            .sr(N__48553));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_11_4  (
            .in0(N__34248),
            .in1(N__30706),
            .in2(_gnd_net_),
            .in3(N__30689),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49082),
            .ce(),
            .sr(N__48553));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_11_5  (
            .in0(N__34191),
            .in1(N__30676),
            .in2(_gnd_net_),
            .in3(N__30662),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49082),
            .ce(),
            .sr(N__48553));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_11_6  (
            .in0(N__34249),
            .in1(N__30657),
            .in2(_gnd_net_),
            .in3(N__30641),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49082),
            .ce(),
            .sr(N__48553));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_11_7  (
            .in0(N__34192),
            .in1(N__30636),
            .in2(_gnd_net_),
            .in3(N__30620),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49082),
            .ce(),
            .sr(N__48553));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_12_0  (
            .in0(N__34200),
            .in1(N__30617),
            .in2(_gnd_net_),
            .in3(N__30599),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49072),
            .ce(),
            .sr(N__48564));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_12_1  (
            .in0(N__34205),
            .in1(N__30588),
            .in2(_gnd_net_),
            .in3(N__30566),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49072),
            .ce(),
            .sr(N__48564));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_12_2  (
            .in0(N__34201),
            .in1(N__30562),
            .in2(_gnd_net_),
            .in3(N__30542),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49072),
            .ce(),
            .sr(N__48564));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_12_3  (
            .in0(N__34206),
            .in1(N__30534),
            .in2(_gnd_net_),
            .in3(N__30518),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49072),
            .ce(),
            .sr(N__48564));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_12_4  (
            .in0(N__34202),
            .in1(N__30930),
            .in2(_gnd_net_),
            .in3(N__30914),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49072),
            .ce(),
            .sr(N__48564));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_12_5  (
            .in0(N__34207),
            .in1(N__30905),
            .in2(_gnd_net_),
            .in3(N__30887),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49072),
            .ce(),
            .sr(N__48564));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_12_6  (
            .in0(N__34203),
            .in1(N__30878),
            .in2(_gnd_net_),
            .in3(N__30884),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49072),
            .ce(),
            .sr(N__48564));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_12_7 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_12_7  (
            .in0(N__34943),
            .in1(N__30860),
            .in2(N__30835),
            .in3(N__34204),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49072),
            .ce(),
            .sr(N__48564));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__30845),
            .in2(N__30809),
            .in3(N__30825),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__30800),
            .in2(N__30779),
            .in3(N__30794),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_13_2  (
            .in0(N__30770),
            .in1(N__30752),
            .in2(N__30746),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__30713),
            .in2(N__30737),
            .in3(N__30728),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_13_4  (
            .in0(N__31187),
            .in1(N__31172),
            .in2(N__31157),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_13_5  (
            .in0(N__31148),
            .in1(N__31133),
            .in2(N__31121),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__31112),
            .in2(N__31082),
            .in3(N__31100),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__31073),
            .in2(N__31043),
            .in3(N__31061),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__31031),
            .in2(N__31004),
            .in3(N__31019),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__32609),
            .in2(N__30980),
            .in3(N__30995),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__30971),
            .in2(N__30941),
            .in3(N__30956),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__31364),
            .in2(N__31394),
            .in3(N__31379),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_14_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_14_4  (
            .in0(N__31358),
            .in1(N__31343),
            .in2(N__31331),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_14_5  (
            .in0(N__31319),
            .in1(N__32822),
            .in2(N__31304),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_14_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_14_6  (
            .in0(N__31295),
            .in1(N__31280),
            .in2(N__31271),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__32597),
            .in2(N__32525),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__31262),
            .in2(N__31250),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__31232),
            .in2(N__31223),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__31208),
            .in2(N__31199),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__31622),
            .in2(N__31613),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__31601),
            .in2(N__31592),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__31574),
            .in2(N__31562),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_11_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_11_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__31547),
            .in2(N__31535),
            .in3(N__31499),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31496),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_11_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_11_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__31489),
            .in2(_gnd_net_),
            .in3(N__35233),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_11_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_11_16_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_11_16_1  (
            .in0(N__35231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31465),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_16_2  (
            .in0(N__31440),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35238),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_16_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_16_3  (
            .in0(N__35236),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31414),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_11_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_11_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_11_16_4  (
            .in0(N__32503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35237),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_16_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_16_5  (
            .in0(N__35234),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32479),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_11_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_11_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_11_16_6  (
            .in0(N__32455),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35232),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_11_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_11_16_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_11_16_7  (
            .in0(N__35235),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32428),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_11_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_11_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_11_17_2 .LUT_INIT=16'b0100010001010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_11_17_2  (
            .in0(N__32408),
            .in1(N__32384),
            .in2(N__32225),
            .in3(N__32031),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49038),
            .ce(),
            .sr(N__48609));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_11_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_11_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33481),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49038),
            .ce(),
            .sr(N__48609));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_11_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_11_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_11_17_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_11_17_7  (
            .in0(N__35253),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49038),
            .ce(),
            .sr(N__48609));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_18_6  (
            .in0(N__31691),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31658),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_4_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_4_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_12_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32741),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49128),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_12_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_12_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_12_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_22_LC_12_7_5  (
            .in0(N__32730),
            .in1(N__32708),
            .in2(_gnd_net_),
            .in3(N__34586),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49106),
            .ce(N__34184),
            .sr(N__48525));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_12_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_12_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_12_8_0  (
            .in0(N__34625),
            .in1(N__32662),
            .in2(_gnd_net_),
            .in3(N__32638),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_8_4  (
            .in0(N__34624),
            .in1(N__34767),
            .in2(_gnd_net_),
            .in3(N__34743),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_12_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_12_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_12_9_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_12_9_1  (
            .in0(N__32883),
            .in1(_gnd_net_),
            .in2(N__32930),
            .in3(N__34683),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49089),
            .ce(N__34185),
            .sr(N__48534));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_12_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_12_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_12_9_2  (
            .in0(N__34681),
            .in1(N__32769),
            .in2(_gnd_net_),
            .in3(N__32809),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49089),
            .ce(N__34185),
            .sr(N__48534));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_12_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_12_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_12_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_12_9_7  (
            .in0(N__32658),
            .in1(N__32642),
            .in2(_gnd_net_),
            .in3(N__34682),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49089),
            .ce(N__34185),
            .sr(N__48534));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_0  (
            .in0(N__32562),
            .in1(N__32537),
            .in2(N__32585),
            .in3(N__32548),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_10_1 .LUT_INIT=16'b1111011101010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_10_1  (
            .in0(N__32580),
            .in1(N__32563),
            .in2(N__32549),
            .in3(N__32536),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_10_2  (
            .in0(N__34612),
            .in1(N__32887),
            .in2(_gnd_net_),
            .in3(N__32929),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_10_3  (
            .in0(N__32848),
            .in1(N__34613),
            .in2(_gnd_net_),
            .in3(N__32866),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_12_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_12_10_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__34611),
            .in2(N__32852),
            .in3(N__32849),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49080),
            .ce(N__34258),
            .sr(N__48541));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_10_6  (
            .in0(N__32810),
            .in1(N__34610),
            .in2(_gnd_net_),
            .in3(N__32773),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__33731),
            .in2(N__33692),
            .in3(N__33690),
            .lcout(\current_shift_inst.control_input_18 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__33803),
            .in2(_gnd_net_),
            .in3(N__32753),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__33797),
            .in2(_gnd_net_),
            .in3(N__32750),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__33791),
            .in2(_gnd_net_),
            .in3(N__32747),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__33785),
            .in2(_gnd_net_),
            .in3(N__32744),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__33779),
            .in2(_gnd_net_),
            .in3(N__32957),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__33773),
            .in2(_gnd_net_),
            .in3(N__32954),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__33767),
            .in2(_gnd_net_),
            .in3(N__32951),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__33761),
            .in2(_gnd_net_),
            .in3(N__32948),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__33755),
            .in2(_gnd_net_),
            .in3(N__32945),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__33122),
            .in2(_gnd_net_),
            .in3(N__32942),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__36161),
            .in2(_gnd_net_),
            .in3(N__32939),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__33671),
            .in2(_gnd_net_),
            .in3(N__32936),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__44471),
            .in2(_gnd_net_),
            .in3(N__32933),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_12_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_12_7  (
            .in0(N__36098),
            .in1(N__36191),
            .in2(_gnd_net_),
            .in3(N__44470),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__33107),
            .in2(_gnd_net_),
            .in3(N__33116),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__33101),
            .in2(_gnd_net_),
            .in3(N__33071),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__49060),
            .ce(),
            .sr(N__48565));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_13_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33068),
            .in3(N__33035),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__49060),
            .ce(),
            .sr(N__48565));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__33032),
            .in2(_gnd_net_),
            .in3(N__33023),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__49060),
            .ce(),
            .sr(N__48565));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__33020),
            .in2(_gnd_net_),
            .in3(N__32984),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__49060),
            .ce(),
            .sr(N__48565));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__32981),
            .in2(_gnd_net_),
            .in3(N__32972),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__49060),
            .ce(),
            .sr(N__48565));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__32969),
            .in2(_gnd_net_),
            .in3(N__32960),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__49060),
            .ce(),
            .sr(N__48565));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__33257),
            .in2(_gnd_net_),
            .in3(N__33248),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__49060),
            .ce(),
            .sr(N__48565));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__33245),
            .in2(_gnd_net_),
            .in3(N__33236),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__49052),
            .ce(),
            .sr(N__48574));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__33233),
            .in2(_gnd_net_),
            .in3(N__33224),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__49052),
            .ce(),
            .sr(N__48574));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__33221),
            .in2(_gnd_net_),
            .in3(N__33212),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__49052),
            .ce(),
            .sr(N__48574));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__33209),
            .in2(_gnd_net_),
            .in3(N__33200),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__49052),
            .ce(),
            .sr(N__48574));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__33197),
            .in2(_gnd_net_),
            .in3(N__33164),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__49052),
            .ce(),
            .sr(N__48574));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_12_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_12_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_12_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__33971),
            .in2(_gnd_net_),
            .in3(N__33161),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__49052),
            .ce(),
            .sr(N__48574));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_12_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_12_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_12_14_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__33986),
            .in2(_gnd_net_),
            .in3(N__33158),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49052),
            .ce(),
            .sr(N__48574));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_12_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_12_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_12_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33151),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49052),
            .ce(),
            .sr(N__48574));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33507),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33465),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_12_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_12_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_12_15_2  (
            .in0(N__35176),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33432),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_12_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_12_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__33405),
            .in2(_gnd_net_),
            .in3(N__35177),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33372),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_15_5  (
            .in0(N__33342),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35174),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_15_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_15_6  (
            .in0(N__35175),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33318),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_12_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_12_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33282),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_12_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_12_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_12_16_0 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst1.state_0_LC_12_16_0  (
            .in0(N__35881),
            .in1(N__34903),
            .in2(N__34888),
            .in3(N__33565),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49037),
            .ce(),
            .sr(N__48590));
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_12_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_12_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a2_1_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__35058),
            .in2(_gnd_net_),
            .in3(N__34818),
            .lcout(state_ns_i_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__34902),
            .in2(_gnd_net_),
            .in3(N__33564),
            .lcout(\phase_controller_inst1.N_55 ),
            .ltout(\phase_controller_inst1.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_12_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_12_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_12_16_3 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \phase_controller_inst1.state_3_LC_12_16_3  (
            .in0(N__36336),
            .in1(N__39219),
            .in2(N__33662),
            .in3(N__33652),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49037),
            .ce(),
            .sr(N__48590));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_17_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__35239),
            .in2(_gnd_net_),
            .in3(N__33636),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_17_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_17_4  (
            .in0(N__36337),
            .in1(N__39195),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_1_LC_12_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_12_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_12_18_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \phase_controller_inst1.state_1_LC_12_18_0  (
            .in0(N__34796),
            .in1(N__34884),
            .in2(_gnd_net_),
            .in3(N__35872),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49026),
            .ce(),
            .sr(N__48610));
    defparam \phase_controller_inst2.start_timer_hc_LC_12_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_12_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_12_18_5 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_12_18_5  (
            .in0(N__34837),
            .in1(N__33617),
            .in2(N__35804),
            .in3(N__33602),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49026),
            .ce(),
            .sr(N__48610));
    defparam \phase_controller_inst1.T23_LC_12_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.T23_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T23_LC_12_19_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst1.T23_LC_12_19_1  (
            .in0(N__33583),
            .in1(N__35873),
            .in2(_gnd_net_),
            .in3(N__33571),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49021),
            .ce(),
            .sr(N__48618));
    defparam \phase_controller_inst1.T45_LC_12_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.T45_LC_12_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T45_LC_12_19_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \phase_controller_inst1.T45_LC_12_19_6  (
            .in0(N__33572),
            .in1(N__33535),
            .in2(_gnd_net_),
            .in3(N__39214),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49021),
            .ce(),
            .sr(N__48618));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_21_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_21_0  (
            .in0(N__41023),
            .in1(N__40986),
            .in2(_gnd_net_),
            .in3(N__49336),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_25_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_25_6  (
            .in0(_gnd_net_),
            .in1(N__37049),
            .in2(_gnd_net_),
            .in3(N__35811),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_26_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_26_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_12_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35813),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49008),
            .ce(),
            .sr(N__48656));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_6_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__34975),
            .in2(_gnd_net_),
            .in3(N__35092),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_8_0 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_8_0  (
            .in0(N__42165),
            .in1(N__44305),
            .in2(N__41411),
            .in3(N__44728),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_8_1 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_8_1  (
            .in0(N__44733),
            .in1(N__46646),
            .in2(N__41705),
            .in3(N__42163),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_8_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_8_2  (
            .in0(N__42161),
            .in1(N__44735),
            .in2(N__46328),
            .in3(N__39110),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_8_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_8_3  (
            .in0(N__44729),
            .in1(N__42166),
            .in2(N__44234),
            .in3(N__41542),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_8_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_8_4  (
            .in0(N__45694),
            .in1(N__44730),
            .in2(N__42319),
            .in3(N__41332),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_8_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_8_5  (
            .in0(N__44732),
            .in1(N__42162),
            .in2(N__46724),
            .in3(N__38980),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_8_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_8_6  (
            .in0(N__42164),
            .in1(N__44731),
            .in2(N__41582),
            .in3(N__45170),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_8_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_8_7  (
            .in0(N__44734),
            .in1(N__46574),
            .in2(N__42320),
            .in3(N__38948),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_13_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_13_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_13_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33965),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49100),
            .ce(),
            .sr(N__48529));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_10_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_10_0  (
            .in0(N__45479),
            .in1(N__41864),
            .in2(_gnd_net_),
            .in3(N__38911),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45478),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_10_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_10_2  (
            .in0(N__35912),
            .in1(N__36152),
            .in2(_gnd_net_),
            .in3(N__44426),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_13_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_13_10_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33725),
            .in3(N__33691),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49092),
            .ce(),
            .sr(N__48535));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_13_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_13_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44427),
            .lcout(\current_shift_inst.N_1326_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44429),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_10_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_10_7  (
            .in0(N__44428),
            .in1(N__36143),
            .in2(_gnd_net_),
            .in3(N__35897),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_11_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_11_0  (
            .in0(N__36134),
            .in1(N__36050),
            .in2(_gnd_net_),
            .in3(N__44462),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_11_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_11_1  (
            .in0(N__44463),
            .in1(N__36125),
            .in2(_gnd_net_),
            .in3(N__36035),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_11_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_11_2  (
            .in0(N__36011),
            .in1(N__36116),
            .in2(_gnd_net_),
            .in3(N__44464),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_11_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_11_3  (
            .in0(N__44465),
            .in1(N__35990),
            .in2(_gnd_net_),
            .in3(N__36236),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_11_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_11_4  (
            .in0(N__35966),
            .in1(N__36227),
            .in2(_gnd_net_),
            .in3(N__44466),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_11_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_11_5  (
            .in0(N__44467),
            .in1(N__35954),
            .in2(_gnd_net_),
            .in3(N__36218),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_11_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_11_6  (
            .in0(N__35942),
            .in1(N__36209),
            .in2(_gnd_net_),
            .in3(N__44468),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_11_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_11_7  (
            .in0(N__44469),
            .in1(N__35924),
            .in2(_gnd_net_),
            .in3(N__36200),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_13_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_13_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_21_LC_13_12_7  (
            .in0(N__34772),
            .in1(N__34745),
            .in2(_gnd_net_),
            .in3(N__34687),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49073),
            .ce(N__34155),
            .sr(N__48546));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_13_13_0  (
            .in0(N__49452),
            .in1(N__35768),
            .in2(_gnd_net_),
            .in3(N__40214),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49066),
            .ce(N__49982),
            .sr(N__48554));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_1  (
            .in0(N__36300),
            .in1(N__39932),
            .in2(_gnd_net_),
            .in3(N__49453),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49066),
            .ce(N__49982),
            .sr(N__48554));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33982),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33951),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33912),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33867),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35651),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33825),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_14_6  (
            .in0(N__35121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35217),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_LC_13_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_15_1 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_13_15_1  (
            .in0(N__34820),
            .in1(N__35105),
            .in2(N__34850),
            .in3(N__35088),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49053),
            .ce(),
            .sr(N__48575));
    defparam \phase_controller_inst1.state_4_LC_13_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_13_15_4 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_13_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__35037),
            .in2(_gnd_net_),
            .in3(N__34819),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49053),
            .ce(),
            .sr(N__48575));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7 .LUT_INIT=16'b1101000011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7  (
            .in0(N__35002),
            .in1(N__34904),
            .in2(N__34982),
            .in3(N__34942),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49053),
            .ce(),
            .sr(N__48575));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_16_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_16_0  (
            .in0(N__35880),
            .in1(N__39167),
            .in2(N__34889),
            .in3(N__39253),
            .lcout(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_13_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_13_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_13_16_1  (
            .in0(N__39279),
            .in1(N__40279),
            .in2(_gnd_net_),
            .in3(N__49429),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_13_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_13_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__39166),
            .in2(_gnd_net_),
            .in3(N__39252),
            .lcout(\phase_controller_inst1.N_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_13_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_17_4 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_13_17_4  (
            .in0(N__34836),
            .in1(N__34792),
            .in2(N__34781),
            .in3(N__50132),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49039),
            .ce(),
            .sr(N__48591));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50133),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49039),
            .ce(),
            .sr(N__48591));
    defparam \phase_controller_inst1.T12_LC_13_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.T12_LC_13_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T12_LC_13_17_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst1.T12_LC_13_17_7  (
            .in0(N__35494),
            .in1(N__35871),
            .in2(_gnd_net_),
            .in3(N__39172),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49039),
            .ce(),
            .sr(N__48591));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_13_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_13_18_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_13_18_4  (
            .in0(N__36259),
            .in1(N__40075),
            .in2(_gnd_net_),
            .in3(N__49546),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_13_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_13_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_13_18_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_13_18_6  (
            .in0(N__35573),
            .in1(N__40144),
            .in2(_gnd_net_),
            .in3(N__49547),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49031),
            .ce(N__50031),
            .sr(N__48601));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_19_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__40211),
            .in2(_gnd_net_),
            .in3(N__40278),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_19_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_19_1  (
            .in0(N__47095),
            .in1(N__49709),
            .in2(N__35483),
            .in3(N__35480),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_19_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_19_4  (
            .in0(N__43874),
            .in1(N__49418),
            .in2(_gnd_net_),
            .in3(N__40908),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_5 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_5  (
            .in0(N__35650),
            .in1(N__35702),
            .in2(_gnd_net_),
            .in3(N__35680),
            .lcout(\current_shift_inst.timer_s1.N_168_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_19_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_19_6  (
            .in0(N__40001),
            .in1(N__40074),
            .in2(N__39920),
            .in3(N__40139),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_13_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_13_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35472),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_20_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_20_0  (
            .in0(N__35540),
            .in1(N__35549),
            .in2(N__36491),
            .in3(N__36468),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_20_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_20_1  (
            .in0(N__35548),
            .in1(N__36489),
            .in2(N__36470),
            .in3(N__35539),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_13_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_13_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_13_20_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_22_LC_13_20_2  (
            .in0(N__49419),
            .in1(N__43499),
            .in2(_gnd_net_),
            .in3(N__39830),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49022),
            .ce(N__48719),
            .sr(N__48619));
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_13_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_13_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_13_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_23_LC_13_20_3  (
            .in0(N__43529),
            .in1(N__39860),
            .in2(_gnd_net_),
            .in3(N__49421),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49022),
            .ce(N__48719),
            .sr(N__48619));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_13_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_13_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_13_20_7  (
            .in0(N__40070),
            .in1(N__36260),
            .in2(_gnd_net_),
            .in3(N__49420),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49022),
            .ce(N__48719),
            .sr(N__48619));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_21_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_21_0  (
            .in0(N__36405),
            .in1(N__36510),
            .in2(N__35522),
            .in3(N__35531),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_21_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_21_1  (
            .in0(N__35530),
            .in1(N__36406),
            .in2(N__36512),
            .in3(N__35518),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_13_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_13_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_13_21_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_20_LC_13_21_2  (
            .in0(N__48112),
            .in1(N__47595),
            .in2(_gnd_net_),
            .in3(N__49353),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49018),
            .ce(N__48717),
            .sr(N__48626));
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_13_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_13_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_13_21_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_21_LC_13_21_3  (
            .in0(N__47703),
            .in1(N__49350),
            .in2(_gnd_net_),
            .in3(N__47686),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49018),
            .ce(N__48717),
            .sr(N__48626));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_13_22_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_13_22_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_13_22_0  (
            .in0(N__49320),
            .in1(N__35568),
            .in2(_gnd_net_),
            .in3(N__40140),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_22_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_22_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_22_1  (
            .in0(N__47599),
            .in1(N__48107),
            .in2(_gnd_net_),
            .in3(N__49318),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_22_2 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_22_2  (
            .in0(N__38309),
            .in1(N__35594),
            .in2(N__48023),
            .in3(N__41016),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_13_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_13_22_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_13_22_3  (
            .in0(N__47707),
            .in1(_gnd_net_),
            .in2(N__35585),
            .in3(N__47679),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_22_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_22_5  (
            .in0(N__50197),
            .in1(N__50172),
            .in2(_gnd_net_),
            .in3(N__49321),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_22_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_22_6  (
            .in0(N__49319),
            .in1(N__35763),
            .in2(_gnd_net_),
            .in3(N__40212),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_13_23_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_13_23_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_13_23_2  (
            .in0(N__43840),
            .in1(N__49335),
            .in2(_gnd_net_),
            .in3(N__47809),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(N__35646),
            .in2(_gnd_net_),
            .in3(N__35679),
            .lcout(\current_shift_inst.timer_s1.N_167_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_23_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_23_4  (
            .in0(N__36280),
            .in1(N__40002),
            .in2(_gnd_net_),
            .in3(N__49334),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_13_24_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_13_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_13_24_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_13_24_0  (
            .in0(N__49573),
            .in1(N__35569),
            .in2(_gnd_net_),
            .in3(N__40145),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49012),
            .ce(N__48712),
            .sr(N__48642));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_13_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_13_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_13_24_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_13_24_1  (
            .in0(N__39280),
            .in1(_gnd_net_),
            .in2(N__49578),
            .in3(N__40280),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49012),
            .ce(N__48712),
            .sr(N__48642));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_13_24_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_13_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_13_24_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_13_24_3  (
            .in0(N__35764),
            .in1(_gnd_net_),
            .in2(N__49579),
            .in3(N__40213),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49012),
            .ce(N__48712),
            .sr(N__48642));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_13_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_13_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_13_24_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_13_24_4  (
            .in0(N__49572),
            .in1(N__43836),
            .in2(_gnd_net_),
            .in3(N__47810),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49012),
            .ce(N__48712),
            .sr(N__48642));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_13_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_13_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_13_24_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_13_24_5  (
            .in0(N__49469),
            .in1(N__36276),
            .in2(_gnd_net_),
            .in3(N__40003),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49012),
            .ce(N__48712),
            .sr(N__48642));
    defparam \current_shift_inst.stop_timer_s1_LC_13_25_2 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_13_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_13_25_2 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_13_25_2  (
            .in0(N__35608),
            .in1(N__39229),
            .in2(N__35681),
            .in3(N__35700),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49011),
            .ce(),
            .sr(N__48647));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_13_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_13_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_13_25_3 .LUT_INIT=16'b1101110000001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_13_25_3  (
            .in0(N__37067),
            .in1(N__35724),
            .in2(N__37277),
            .in3(N__37051),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49011),
            .ce(),
            .sr(N__48647));
    defparam \current_shift_inst.start_timer_s1_LC_13_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_13_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_13_25_4 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_13_25_4  (
            .in0(N__35607),
            .in1(N__35699),
            .in2(_gnd_net_),
            .in3(N__39228),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49011),
            .ce(),
            .sr(N__48647));
    defparam \current_shift_inst.timer_s1.running_LC_13_25_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_25_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_25_5  (
            .in0(N__35701),
            .in1(N__35675),
            .in2(_gnd_net_),
            .in3(N__35645),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49011),
            .ce(),
            .sr(N__48647));
    defparam \phase_controller_inst1.S1_LC_13_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_13_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39230),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49011),
            .ce(),
            .sr(N__48647));
    defparam \phase_controller_inst2.stoper_hc.running_LC_13_26_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_13_26_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_13_26_1 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_13_26_1  (
            .in0(N__37050),
            .in1(N__37066),
            .in2(N__35828),
            .in3(N__37273),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49009),
            .ce(),
            .sr(N__48650));
    defparam \phase_controller_inst1.S2_LC_13_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_26_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35885),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49009),
            .ce(),
            .sr(N__48650));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_27_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_27_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_27_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_27_5  (
            .in0(N__37048),
            .in1(N__35824),
            .in2(_gnd_net_),
            .in3(N__35812),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_13_27_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_13_27_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_13_27_7 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_13_27_7  (
            .in0(N__38553),
            .in1(N__40889),
            .in2(N__38600),
            .in3(N__40959),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_4_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_4_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_14_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39594),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35777),
            .ce(),
            .sr(N__48517));
    defparam \delay_measurement_inst.start_timer_hc_LC_14_4_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_14_4_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_14_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_14_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39593),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35777),
            .ce(),
            .sr(N__48517));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_5_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(N__37622),
            .in2(N__37640),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_5_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__37590),
            .in2(N__37205),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_5_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__42213),
            .in2(N__37496),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_5_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(N__37523),
            .in2(N__42387),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_5_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(N__42217),
            .in2(N__37217),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_5_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(N__37544),
            .in2(N__42388),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_5_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(N__42221),
            .in2(N__37178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_5_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__37550),
            .in2(N__42389),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_6_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(N__42225),
            .in2(N__37187),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_6_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__37166),
            .in2(N__42390),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_6_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__42229),
            .in2(N__37532),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_6_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__38771),
            .in2(N__42391),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_6_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__42233),
            .in2(N__38762),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_6_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__38483),
            .in2(N__42392),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_6_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(N__42237),
            .in2(N__37196),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_6_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__38492),
            .in2(N__42393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_7_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__42241),
            .in2(N__38726),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_7_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__42245),
            .in2(N__37706),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_7_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__42242),
            .in2(N__38714),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_7_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__42246),
            .in2(N__39047),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_7_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__42243),
            .in2(N__38750),
            .in3(N__35900),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_7_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__42247),
            .in2(N__41894),
            .in3(N__35888),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_7_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__42244),
            .in2(N__38738),
            .in3(N__36038),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_7_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__42248),
            .in2(N__38699),
            .in3(N__36023),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__42131),
            .in2(N__36020),
            .in3(N__35999),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__35996),
            .in2(N__42303),
            .in3(N__35978),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__42135),
            .in2(N__35975),
            .in3(N__35957),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__37517),
            .in2(N__42304),
            .in3(N__35945),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__42139),
            .in2(N__42530),
            .in3(N__35933),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__35930),
            .in2(N__42305),
            .in3(N__35915),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__42143),
            .in2(N__37724),
            .in3(N__36086),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_8_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_8_7  (
            .in0(N__42144),
            .in1(N__44752),
            .in2(_gnd_net_),
            .in3(N__36083),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__37615),
            .in2(N__37484),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_9_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_9_1  (
            .in0(N__43798),
            .in1(N__37583),
            .in2(N__37559),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__42103),
            .in2(N__37508),
            .in3(N__43799),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__36080),
            .in2(N__42296),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__42107),
            .in2(N__36068),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__38504),
            .in2(N__42297),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__42111),
            .in2(N__36059),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__40844),
            .in2(N__42298),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__42115),
            .in2(N__37685),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__37781),
            .in2(N__42299),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__42119),
            .in2(N__37793),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__37775),
            .in2(N__42300),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(N__42123),
            .in2(N__37715),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__36107),
            .in2(N__42301),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(N__42127),
            .in2(N__37694),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__37730),
            .in2(N__42302),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__42249),
            .in2(N__37811),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__37754),
            .in2(N__42394),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(N__42253),
            .in2(N__37748),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__37769),
            .in2(N__42395),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__42257),
            .in2(N__37739),
            .in3(N__36146),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__42485),
            .in2(N__42396),
            .in3(N__36137),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(N__42261),
            .in2(N__37763),
            .in3(N__36128),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__39056),
            .in2(N__42397),
            .in3(N__36119),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__42306),
            .in2(N__37850),
            .in3(N__36110),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__37835),
            .in2(N__42422),
            .in3(N__36230),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__42310),
            .in2(N__37829),
            .in3(N__36221),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__37802),
            .in2(N__42423),
            .in3(N__36212),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__42314),
            .in2(N__37862),
            .in3(N__36203),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__37841),
            .in2(N__42424),
            .in3(N__36194),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__42318),
            .in2(N__37820),
            .in3(N__36182),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_12_7 .LUT_INIT=16'b1000101101000111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_12_7  (
            .in0(N__42497),
            .in1(N__44461),
            .in2(N__36179),
            .in3(N__36164),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_14_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_14_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_14_13_3  (
            .in0(N__36304),
            .in1(N__39928),
            .in2(_gnd_net_),
            .in3(N__49580),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_14_14_7 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_14_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48680),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_2_LC_14_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_14_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_14_16_6 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_14_16_6  (
            .in0(N__39215),
            .in1(N__39168),
            .in2(N__36341),
            .in3(N__39254),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49054),
            .ce(),
            .sr(N__48576));
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_14_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_14_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_24_LC_14_17_2  (
            .in0(N__49479),
            .in1(N__47378),
            .in2(_gnd_net_),
            .in3(N__47396),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49047),
            .ce(N__48722),
            .sr(N__48584));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_14_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_14_17_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_14_17_3  (
            .in0(N__36308),
            .in1(N__39927),
            .in2(_gnd_net_),
            .in3(N__49481),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49047),
            .ce(N__48722),
            .sr(N__48584));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_14_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_14_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_14_17_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_14_17_7  (
            .in0(N__47850),
            .in1(N__49480),
            .in2(_gnd_net_),
            .in3(N__46913),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49047),
            .ce(N__48722),
            .sr(N__48584));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_14_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_14_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_14_18_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_14_18_1  (
            .in0(N__36284),
            .in1(N__40004),
            .in2(_gnd_net_),
            .in3(N__49550),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49040),
            .ce(N__50027),
            .sr(N__48592));
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_14_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_14_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_14_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_31_LC_14_18_2  (
            .in0(N__49548),
            .in1(N__41027),
            .in2(_gnd_net_),
            .in3(N__40990),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49040),
            .ce(N__50027),
            .sr(N__48592));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_14_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_14_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_14_18_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_14_18_5  (
            .in0(N__36255),
            .in1(N__40076),
            .in2(_gnd_net_),
            .in3(N__49549),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49040),
            .ce(N__50027),
            .sr(N__48592));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__37247),
            .in2(N__37466),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_19_1  (
            .in0(N__37417),
            .in1(N__36538),
            .in2(_gnd_net_),
            .in3(N__36239),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49032),
            .ce(),
            .sr(N__48602));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_19_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_19_2  (
            .in0(N__37425),
            .in1(N__36805),
            .in2(N__37454),
            .in3(N__36389),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49032),
            .ce(),
            .sr(N__48602));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_19_3  (
            .in0(N__37418),
            .in1(N__36781),
            .in2(_gnd_net_),
            .in3(N__36386),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49032),
            .ce(),
            .sr(N__48602));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_19_4  (
            .in0(N__37426),
            .in1(N__36754),
            .in2(_gnd_net_),
            .in3(N__36383),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49032),
            .ce(),
            .sr(N__48602));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_19_5  (
            .in0(N__37419),
            .in1(N__36730),
            .in2(_gnd_net_),
            .in3(N__36380),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49032),
            .ce(),
            .sr(N__48602));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_19_6  (
            .in0(N__37427),
            .in1(N__36700),
            .in2(_gnd_net_),
            .in3(N__36377),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49032),
            .ce(),
            .sr(N__48602));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_19_7  (
            .in0(N__37420),
            .in1(N__36670),
            .in2(_gnd_net_),
            .in3(N__36374),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49032),
            .ce(),
            .sr(N__48602));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_20_0  (
            .in0(N__37431),
            .in1(N__36640),
            .in2(_gnd_net_),
            .in3(N__36371),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49027),
            .ce(),
            .sr(N__48611));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_20_1  (
            .in0(N__37413),
            .in1(N__37003),
            .in2(_gnd_net_),
            .in3(N__36368),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49027),
            .ce(),
            .sr(N__48611));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_20_2  (
            .in0(N__37428),
            .in1(N__36961),
            .in2(_gnd_net_),
            .in3(N__36365),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49027),
            .ce(),
            .sr(N__48611));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_20_3  (
            .in0(N__37414),
            .in1(N__36925),
            .in2(_gnd_net_),
            .in3(N__36431),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49027),
            .ce(),
            .sr(N__48611));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_20_4  (
            .in0(N__37429),
            .in1(N__36892),
            .in2(_gnd_net_),
            .in3(N__36428),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49027),
            .ce(),
            .sr(N__48611));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_20_5  (
            .in0(N__37415),
            .in1(N__36856),
            .in2(_gnd_net_),
            .in3(N__36425),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49027),
            .ce(),
            .sr(N__48611));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_20_6  (
            .in0(N__37430),
            .in1(N__36829),
            .in2(_gnd_net_),
            .in3(N__36422),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49027),
            .ce(),
            .sr(N__48611));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_20_7  (
            .in0(N__37416),
            .in1(N__38261),
            .in2(_gnd_net_),
            .in3(N__36419),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49027),
            .ce(),
            .sr(N__48611));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_21_0  (
            .in0(N__37421),
            .in1(N__38241),
            .in2(_gnd_net_),
            .in3(N__36416),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49023),
            .ce(),
            .sr(N__48620));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_21_1  (
            .in0(N__37432),
            .in1(N__38665),
            .in2(_gnd_net_),
            .in3(N__36413),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49023),
            .ce(),
            .sr(N__48620));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_21_2  (
            .in0(N__37422),
            .in1(N__38641),
            .in2(_gnd_net_),
            .in3(N__36410),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49023),
            .ce(),
            .sr(N__48620));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_21_3  (
            .in0(N__37433),
            .in1(N__36407),
            .in2(_gnd_net_),
            .in3(N__36392),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49023),
            .ce(),
            .sr(N__48620));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_21_4  (
            .in0(N__37423),
            .in1(N__36511),
            .in2(_gnd_net_),
            .in3(N__36494),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49023),
            .ce(),
            .sr(N__48620));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_21_5  (
            .in0(N__37434),
            .in1(N__36490),
            .in2(_gnd_net_),
            .in3(N__36473),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49023),
            .ce(),
            .sr(N__48620));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_21_6  (
            .in0(N__37424),
            .in1(N__36469),
            .in2(_gnd_net_),
            .in3(N__36452),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49023),
            .ce(),
            .sr(N__48620));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_21_7  (
            .in0(N__37435),
            .in1(N__36579),
            .in2(_gnd_net_),
            .in3(N__36449),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49023),
            .ce(),
            .sr(N__48620));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_22_0  (
            .in0(N__37402),
            .in1(N__36599),
            .in2(_gnd_net_),
            .in3(N__36446),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49019),
            .ce(),
            .sr(N__48627));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_22_1  (
            .in0(N__37406),
            .in1(N__38474),
            .in2(_gnd_net_),
            .in3(N__36443),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49019),
            .ce(),
            .sr(N__48627));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_22_2  (
            .in0(N__37403),
            .in1(N__38451),
            .in2(_gnd_net_),
            .in3(N__36440),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49019),
            .ce(),
            .sr(N__48627));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_22_3  (
            .in0(N__37407),
            .in1(N__38405),
            .in2(_gnd_net_),
            .in3(N__36437),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49019),
            .ce(),
            .sr(N__48627));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_22_4  (
            .in0(N__37404),
            .in1(N__38389),
            .in2(_gnd_net_),
            .in3(N__36434),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49019),
            .ce(),
            .sr(N__48627));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_22_5  (
            .in0(N__37408),
            .in1(N__38543),
            .in2(_gnd_net_),
            .in3(N__36617),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49019),
            .ce(),
            .sr(N__48627));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_22_6  (
            .in0(N__37405),
            .in1(N__38582),
            .in2(_gnd_net_),
            .in3(N__36614),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49019),
            .ce(),
            .sr(N__48627));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_23_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_23_0  (
            .in0(N__36598),
            .in1(N__36580),
            .in2(N__36563),
            .in3(N__36611),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_14_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_14_23_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_14_23_1  (
            .in0(N__36610),
            .in1(N__36597),
            .in2(N__36584),
            .in3(N__36559),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_14_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_14_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_14_23_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_25_LC_14_23_3  (
            .in0(N__47918),
            .in1(N__47959),
            .in2(_gnd_net_),
            .in3(N__49352),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49014),
            .ce(N__48714),
            .sr(N__48633));
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_14_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_14_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_14_23_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_26_LC_14_23_6  (
            .in0(N__49351),
            .in1(N__50193),
            .in2(_gnd_net_),
            .in3(N__50177),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49014),
            .ce(N__48714),
            .sr(N__48633));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_14_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_14_23_7 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_14_23_7  (
            .in0(N__38299),
            .in1(N__38473),
            .in2(N__38455),
            .in3(N__38341),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_14_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_14_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_14_24_0  (
            .in0(_gnd_net_),
            .in1(N__38324),
            .in2(N__36551),
            .in3(N__37243),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_14_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_14_24_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_14_24_1  (
            .in0(N__36542),
            .in1(N__38612),
            .in2(N__36524),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_14_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_14_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_14_24_2  (
            .in0(_gnd_net_),
            .in1(N__36791),
            .in2(N__38351),
            .in3(N__36809),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_14_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_14_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(N__38330),
            .in2(N__36767),
            .in3(N__36785),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_14_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_14_24_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_14_24_4  (
            .in0(_gnd_net_),
            .in1(N__49157),
            .in2(N__36740),
            .in3(N__36758),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_14_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_14_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(N__38357),
            .in2(N__36716),
            .in3(N__36731),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_14_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_14_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_14_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_14_24_6  (
            .in0(_gnd_net_),
            .in1(N__36707),
            .in2(N__36686),
            .in3(N__36701),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_14_24_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_14_24_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(N__36677),
            .in2(N__36656),
            .in3(N__36671),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_14_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_14_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(N__36647),
            .in2(N__36626),
            .in3(N__36641),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_14_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_14_25_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_14_25_1  (
            .in0(N__37004),
            .in1(N__36989),
            .in2(N__36977),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_14_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_14_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(N__36968),
            .in2(N__36947),
            .in3(N__36962),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_14_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_14_25_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(N__36911),
            .in2(N__36938),
            .in3(N__36926),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_14_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_14_25_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_14_25_4  (
            .in0(_gnd_net_),
            .in1(N__36878),
            .in2(N__36905),
            .in3(N__36896),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_14_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_14_25_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__36872),
            .in2(N__36842),
            .in3(N__36857),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_14_25_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_14_25_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_14_25_6  (
            .in0(N__36830),
            .in1(N__36815),
            .in2(N__40856),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_14_25_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_14_25_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_14_25_7  (
            .in0(_gnd_net_),
            .in1(N__38273),
            .in2(N__38225),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_14_26_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_14_26_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_14_26_0  (
            .in0(_gnd_net_),
            .in1(N__38618),
            .in2(N__38684),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_14_26_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_14_26_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(N__37160),
            .in2(N__37148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_14_26_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_14_26_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_14_26_2  (
            .in0(_gnd_net_),
            .in1(N__37133),
            .in2(N__37121),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_14_26_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_14_26_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(N__37103),
            .in2(N__37094),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_14_26_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_14_26_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_14_26_4  (
            .in0(_gnd_net_),
            .in1(N__37082),
            .in2(N__38429),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_14_26_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_14_26_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_14_26_5  (
            .in0(_gnd_net_),
            .in1(N__38414),
            .in2(N__38372),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_14_26_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_14_26_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_14_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_14_26_6  (
            .in0(_gnd_net_),
            .in1(N__38606),
            .in2(N__38519),
            .in3(N__37073),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_26_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_26_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37070),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_14_27_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_14_27_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_14_27_1 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_14_27_1  (
            .in0(N__38515),
            .in1(N__37055),
            .in2(N__37019),
            .in3(N__37010),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_27_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_27_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_27_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_14_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37469),
            .in3(N__37268),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_14_27_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_14_27_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_14_27_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_14_27_4  (
            .in0(_gnd_net_),
            .in1(N__37267),
            .in2(_gnd_net_),
            .in3(N__37285),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_27_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_27_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_27_6 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_27_6  (
            .in0(N__37409),
            .in1(N__37286),
            .in2(N__37242),
            .in3(N__37269),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49010),
            .ce(),
            .sr(N__48651));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_5_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_5_4 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_5_4  (
            .in0(N__44678),
            .in1(N__42452),
            .in2(N__41543),
            .in3(N__44230),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_15_5_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_15_5_5 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_15_5_5  (
            .in0(N__41384),
            .in1(N__44677),
            .in2(N__37598),
            .in3(N__41362),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_15_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_15_6_0 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_15_6_0  (
            .in0(N__42438),
            .in1(N__44598),
            .in2(N__41207),
            .in3(N__46252),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_6_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_6_1  (
            .in0(N__44595),
            .in1(N__42443),
            .in2(N__45562),
            .in3(N__41308),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_6_2 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_6_2  (
            .in0(N__42441),
            .in1(N__41333),
            .in2(N__45698),
            .in3(N__44593),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_15_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_15_6_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_15_6_3  (
            .in0(N__44596),
            .in1(N__42444),
            .in2(N__38912),
            .in3(N__45477),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_15_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_15_6_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_15_6_4  (
            .in0(N__42442),
            .in1(N__44594),
            .in2(N__41432),
            .in3(N__45626),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_6_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_6_5  (
            .in0(N__44592),
            .in1(N__42440),
            .in2(N__44155),
            .in3(N__41515),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_6_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_6_6  (
            .in0(N__42437),
            .in1(N__44597),
            .in2(N__45404),
            .in3(N__41753),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_15_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_15_6_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_15_6_7  (
            .in0(N__44591),
            .in1(N__42439),
            .in2(N__44309),
            .in3(N__41407),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_7_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_7_1  (
            .in0(N__42325),
            .in1(N__44556),
            .in2(N__46505),
            .in3(N__41606),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_15_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_15_7_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_15_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47135),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49130),
            .ce(N__47168),
            .sr(N__48518));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_7_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_7_3  (
            .in0(N__42326),
            .in1(N__44552),
            .in2(N__44366),
            .in3(N__41182),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_7_4 .LUT_INIT=16'b1010001110100011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_7_4  (
            .in0(N__41183),
            .in1(N__44362),
            .in2(N__44657),
            .in3(N__42327),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_15_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_15_7_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_15_7_5  (
            .in0(N__37667),
            .in1(N__44551),
            .in2(_gnd_net_),
            .in3(N__37676),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_15_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_15_7_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__38826),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_15_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_15_7_7 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__37666),
            .in2(N__37670),
            .in3(N__44550),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44393),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49123),
            .ce(N__47166),
            .sr(N__48519));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_15_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_15_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37664),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_8_2 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_8_2  (
            .in0(N__37665),
            .in1(_gnd_net_),
            .in2(N__37646),
            .in3(N__41847),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_8_4  (
            .in0(N__44890),
            .in1(N__43765),
            .in2(_gnd_net_),
            .in3(N__37604),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_15_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_15_8_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__44891),
            .in2(N__37643),
            .in3(N__37636),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47134),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49123),
            .ce(N__47166),
            .sr(N__48519));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_8_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_8_7  (
            .in0(N__41848),
            .in1(N__45312),
            .in2(_gnd_net_),
            .in3(N__38871),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_9_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_9_0  (
            .in0(N__44658),
            .in1(N__41380),
            .in2(N__37591),
            .in3(N__41352),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_9_1  (
            .in0(N__44335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49116),
            .ce(N__47163),
            .sr(N__48522));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41351),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_9_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__44659),
            .in2(_gnd_net_),
            .in3(N__39075),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_9_6 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_9_6  (
            .in0(N__44660),
            .in1(N__42160),
            .in2(N__39080),
            .in3(N__43800),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_15_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_15_10_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_15_10_0  (
            .in0(N__42182),
            .in1(N__44665),
            .in2(N__45247),
            .in3(N__41491),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_10_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_10_1  (
            .in0(N__44667),
            .in1(N__46037),
            .in2(N__42323),
            .in3(N__41677),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_10_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_10_2  (
            .in0(N__42183),
            .in1(N__44666),
            .in2(N__46256),
            .in3(N__41203),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_10_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_10_3  (
            .in0(N__44668),
            .in1(N__46320),
            .in2(_gnd_net_),
            .in3(N__39102),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_10_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_10_4  (
            .in0(N__42184),
            .in1(N__44661),
            .in2(N__45563),
            .in3(N__41309),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_10_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_10_5  (
            .in0(N__44663),
            .in1(N__45403),
            .in2(N__42321),
            .in3(N__41749),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_10_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_10_6  (
            .in0(N__45476),
            .in1(N__44662),
            .in2(N__42324),
            .in3(N__38904),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_10_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_10_7  (
            .in0(N__44664),
            .in1(N__45322),
            .in2(N__42322),
            .in3(N__38872),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_11_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_11_0  (
            .in0(N__44713),
            .in1(N__45895),
            .in2(N__42469),
            .in3(N__42548),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_11_1 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_11_1  (
            .in0(N__41468),
            .in1(N__42407),
            .in2(N__46865),
            .in3(N__44715),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_15_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_15_11_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_15_11_2  (
            .in0(N__44711),
            .in1(N__46036),
            .in2(N__42468),
            .in3(N__41678),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_11_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_11_3  (
            .in0(N__45967),
            .in1(N__44712),
            .in2(N__41660),
            .in3(N__42416),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_11_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_11_4  (
            .in0(N__44714),
            .in1(N__45823),
            .in2(N__42467),
            .in3(N__41728),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_11_5 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_11_5  (
            .in0(N__41168),
            .in1(N__44710),
            .in2(N__46193),
            .in3(N__42412),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_11_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_11_6  (
            .in0(N__44717),
            .in1(N__46409),
            .in2(N__42466),
            .in3(N__42514),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_11_7 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_11_7  (
            .in0(N__46720),
            .in1(N__44716),
            .in2(N__38987),
            .in3(N__42411),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_12_1 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_12_1  (
            .in0(N__39106),
            .in1(N__46324),
            .in2(N__42471),
            .in3(N__44723),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_12_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_12_2  (
            .in0(N__44720),
            .in1(N__46645),
            .in2(N__42472),
            .in3(N__41698),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_12_3 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_12_3  (
            .in0(N__42431),
            .in1(N__38941),
            .in2(N__46570),
            .in3(N__44721),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_4 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_4  (
            .in0(N__44724),
            .in1(N__42433),
            .in2(N__39079),
            .in3(N__43807),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_12_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_12_5  (
            .in0(N__46563),
            .in1(N__44719),
            .in2(_gnd_net_),
            .in3(N__38940),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_12_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_12_6  (
            .in0(N__44718),
            .in1(N__42432),
            .in2(N__46111),
            .in3(N__42575),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_12_7 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_12_7  (
            .in0(N__41602),
            .in1(N__46501),
            .in2(N__42470),
            .in3(N__44722),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_15_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_15_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_15_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_15_13_0  (
            .in0(N__38125),
            .in1(N__44385),
            .in2(_gnd_net_),
            .in3(N__37796),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__49083),
            .ce(N__38002),
            .sr(N__48542));
    defparam \current_shift_inst.timer_s1.counter_1_LC_15_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_15_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_15_13_1  (
            .in0(N__38117),
            .in1(N__44328),
            .in2(_gnd_net_),
            .in3(N__37889),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__49083),
            .ce(N__38002),
            .sr(N__48542));
    defparam \current_shift_inst.timer_s1.counter_2_LC_15_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_15_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_15_13_2  (
            .in0(N__38126),
            .in1(N__44248),
            .in2(_gnd_net_),
            .in3(N__37886),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__49083),
            .ce(N__38002),
            .sr(N__48542));
    defparam \current_shift_inst.timer_s1.counter_3_LC_15_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_15_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_15_13_3  (
            .in0(N__38118),
            .in1(N__44170),
            .in2(_gnd_net_),
            .in3(N__37883),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__49083),
            .ce(N__38002),
            .sr(N__48542));
    defparam \current_shift_inst.timer_s1.counter_4_LC_15_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_15_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_15_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_15_13_4  (
            .in0(N__38127),
            .in1(N__45714),
            .in2(_gnd_net_),
            .in3(N__37880),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__49083),
            .ce(N__38002),
            .sr(N__48542));
    defparam \current_shift_inst.timer_s1.counter_5_LC_15_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_15_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_15_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_15_13_5  (
            .in0(N__38119),
            .in1(N__45640),
            .in2(_gnd_net_),
            .in3(N__37877),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__49083),
            .ce(N__38002),
            .sr(N__48542));
    defparam \current_shift_inst.timer_s1.counter_6_LC_15_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_15_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_15_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_15_13_6  (
            .in0(N__38128),
            .in1(N__45577),
            .in2(_gnd_net_),
            .in3(N__37874),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__49083),
            .ce(N__38002),
            .sr(N__48542));
    defparam \current_shift_inst.timer_s1.counter_7_LC_15_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_15_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_15_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_15_13_7  (
            .in0(N__38120),
            .in1(N__45493),
            .in2(_gnd_net_),
            .in3(N__37871),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__49083),
            .ce(N__38002),
            .sr(N__48542));
    defparam \current_shift_inst.timer_s1.counter_8_LC_15_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_15_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_15_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_15_14_0  (
            .in0(N__38124),
            .in1(N__45426),
            .in2(_gnd_net_),
            .in3(N__37868),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__49074),
            .ce(N__38003),
            .sr(N__48547));
    defparam \current_shift_inst.timer_s1.counter_9_LC_15_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_15_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_15_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_15_14_1  (
            .in0(N__38132),
            .in1(N__45345),
            .in2(_gnd_net_),
            .in3(N__37865),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__49074),
            .ce(N__38003),
            .sr(N__48547));
    defparam \current_shift_inst.timer_s1.counter_10_LC_15_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_15_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_15_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_15_14_2  (
            .in0(N__38121),
            .in1(N__45264),
            .in2(_gnd_net_),
            .in3(N__37916),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__49074),
            .ce(N__38003),
            .sr(N__48547));
    defparam \current_shift_inst.timer_s1.counter_11_LC_15_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_15_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_15_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_15_14_3  (
            .in0(N__38129),
            .in1(N__45186),
            .in2(_gnd_net_),
            .in3(N__37913),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__49074),
            .ce(N__38003),
            .sr(N__48547));
    defparam \current_shift_inst.timer_s1.counter_12_LC_15_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_15_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_15_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_15_14_4  (
            .in0(N__38122),
            .in1(N__46272),
            .in2(_gnd_net_),
            .in3(N__37910),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__49074),
            .ce(N__38003),
            .sr(N__48547));
    defparam \current_shift_inst.timer_s1.counter_13_LC_15_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_15_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_15_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_15_14_5  (
            .in0(N__38130),
            .in1(N__46207),
            .in2(_gnd_net_),
            .in3(N__37907),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__49074),
            .ce(N__38003),
            .sr(N__48547));
    defparam \current_shift_inst.timer_s1.counter_14_LC_15_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_15_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_15_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_15_14_6  (
            .in0(N__38123),
            .in1(N__46128),
            .in2(_gnd_net_),
            .in3(N__37904),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__49074),
            .ce(N__38003),
            .sr(N__48547));
    defparam \current_shift_inst.timer_s1.counter_15_LC_15_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_15_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_15_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_15_14_7  (
            .in0(N__38131),
            .in1(N__46051),
            .in2(_gnd_net_),
            .in3(N__37901),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__49074),
            .ce(N__38003),
            .sr(N__48547));
    defparam \current_shift_inst.timer_s1.counter_16_LC_15_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_15_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_15_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_15_15_0  (
            .in0(N__38085),
            .in1(N__45987),
            .in2(_gnd_net_),
            .in3(N__37898),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__49067),
            .ce(N__38001),
            .sr(N__48555));
    defparam \current_shift_inst.timer_s1.counter_17_LC_15_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_15_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_15_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_15_15_1  (
            .in0(N__38095),
            .in1(N__45912),
            .in2(_gnd_net_),
            .in3(N__37895),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__49067),
            .ce(N__38001),
            .sr(N__48555));
    defparam \current_shift_inst.timer_s1.counter_18_LC_15_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_15_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_15_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_15_15_2  (
            .in0(N__38086),
            .in1(N__45843),
            .in2(_gnd_net_),
            .in3(N__37892),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__49067),
            .ce(N__38001),
            .sr(N__48555));
    defparam \current_shift_inst.timer_s1.counter_19_LC_15_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_15_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_15_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_15_15_3  (
            .in0(N__38096),
            .in1(N__45771),
            .in2(_gnd_net_),
            .in3(N__37943),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__49067),
            .ce(N__38001),
            .sr(N__48555));
    defparam \current_shift_inst.timer_s1.counter_20_LC_15_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_15_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_15_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_15_15_4  (
            .in0(N__38087),
            .in1(N__46879),
            .in2(_gnd_net_),
            .in3(N__37940),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__49067),
            .ce(N__38001),
            .sr(N__48555));
    defparam \current_shift_inst.timer_s1.counter_21_LC_15_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_15_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_15_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_15_15_5  (
            .in0(N__38097),
            .in1(N__46810),
            .in2(_gnd_net_),
            .in3(N__37937),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__49067),
            .ce(N__38001),
            .sr(N__48555));
    defparam \current_shift_inst.timer_s1.counter_22_LC_15_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_15_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_15_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_15_15_6  (
            .in0(N__38088),
            .in1(N__46738),
            .in2(_gnd_net_),
            .in3(N__37934),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__49067),
            .ce(N__38001),
            .sr(N__48555));
    defparam \current_shift_inst.timer_s1.counter_23_LC_15_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_15_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_15_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_15_15_7  (
            .in0(N__38098),
            .in1(N__46660),
            .in2(_gnd_net_),
            .in3(N__37931),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__49067),
            .ce(N__38001),
            .sr(N__48555));
    defparam \current_shift_inst.timer_s1.counter_24_LC_15_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_15_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_15_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_15_16_0  (
            .in0(N__38089),
            .in1(N__46590),
            .in2(_gnd_net_),
            .in3(N__37928),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__49061),
            .ce(N__37991),
            .sr(N__48566));
    defparam \current_shift_inst.timer_s1.counter_25_LC_15_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_15_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_15_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_15_16_1  (
            .in0(N__38093),
            .in1(N__46521),
            .in2(_gnd_net_),
            .in3(N__37925),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__49061),
            .ce(N__37991),
            .sr(N__48566));
    defparam \current_shift_inst.timer_s1.counter_26_LC_15_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_15_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_15_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_15_16_2  (
            .in0(N__38090),
            .in1(N__46431),
            .in2(_gnd_net_),
            .in3(N__37922),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__49061),
            .ce(N__37991),
            .sr(N__48566));
    defparam \current_shift_inst.timer_s1.counter_27_LC_15_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_15_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_15_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_15_16_3  (
            .in0(N__38094),
            .in1(N__46344),
            .in2(_gnd_net_),
            .in3(N__37919),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__49061),
            .ce(N__37991),
            .sr(N__48566));
    defparam \current_shift_inst.timer_s1.counter_28_LC_15_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_15_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_15_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_15_16_4  (
            .in0(N__38091),
            .in1(N__46450),
            .in2(_gnd_net_),
            .in3(N__38135),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__49061),
            .ce(N__37991),
            .sr(N__48566));
    defparam \current_shift_inst.timer_s1.counter_29_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_15_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_15_16_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_15_16_5  (
            .in0(N__46369),
            .in1(N__38092),
            .in2(_gnd_net_),
            .in3(N__38006),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49061),
            .ce(N__37991),
            .sr(N__48566));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_17_0  (
            .in0(N__39517),
            .in1(N__39789),
            .in2(_gnd_net_),
            .in3(N__37964),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__49055),
            .ce(N__39569),
            .sr(N__48577));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_17_1  (
            .in0(N__39521),
            .in1(N__39732),
            .in2(_gnd_net_),
            .in3(N__37961),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__49055),
            .ce(N__39569),
            .sr(N__48577));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_17_2  (
            .in0(N__39518),
            .in1(N__40353),
            .in2(_gnd_net_),
            .in3(N__37958),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__49055),
            .ce(N__39569),
            .sr(N__48577));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_17_3  (
            .in0(N__39522),
            .in1(N__40321),
            .in2(_gnd_net_),
            .in3(N__37955),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__49055),
            .ce(N__39569),
            .sr(N__48577));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_17_4  (
            .in0(N__39519),
            .in1(N__40299),
            .in2(_gnd_net_),
            .in3(N__37952),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__49055),
            .ce(N__39569),
            .sr(N__48577));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_17_5  (
            .in0(N__39523),
            .in1(N__40230),
            .in2(_gnd_net_),
            .in3(N__37949),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__49055),
            .ce(N__39569),
            .sr(N__48577));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_17_6  (
            .in0(N__39520),
            .in1(N__40161),
            .in2(_gnd_net_),
            .in3(N__37946),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__49055),
            .ce(N__39569),
            .sr(N__48577));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_17_7  (
            .in0(N__39524),
            .in1(N__40092),
            .in2(_gnd_net_),
            .in3(N__38162),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__49055),
            .ce(N__39569),
            .sr(N__48577));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_18_0  (
            .in0(N__39504),
            .in1(N__40023),
            .in2(_gnd_net_),
            .in3(N__38159),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__49048),
            .ce(N__39574),
            .sr(N__48585));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_18_1  (
            .in0(N__39508),
            .in1(N__39951),
            .in2(_gnd_net_),
            .in3(N__38156),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__49048),
            .ce(N__39574),
            .sr(N__48585));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_18_2  (
            .in0(N__39501),
            .in1(N__40596),
            .in2(_gnd_net_),
            .in3(N__38153),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__49048),
            .ce(N__39574),
            .sr(N__48585));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_18_3  (
            .in0(N__39505),
            .in1(N__40575),
            .in2(_gnd_net_),
            .in3(N__38150),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__49048),
            .ce(N__39574),
            .sr(N__48585));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_18_4  (
            .in0(N__39502),
            .in1(N__40551),
            .in2(_gnd_net_),
            .in3(N__38147),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__49048),
            .ce(N__39574),
            .sr(N__48585));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_18_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_18_5  (
            .in0(N__39506),
            .in1(N__40524),
            .in2(_gnd_net_),
            .in3(N__38144),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__49048),
            .ce(N__39574),
            .sr(N__48585));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_18_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_18_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_18_6  (
            .in0(N__39503),
            .in1(N__40494),
            .in2(_gnd_net_),
            .in3(N__38141),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__49048),
            .ce(N__39574),
            .sr(N__48585));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_18_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_18_7  (
            .in0(N__39507),
            .in1(N__40467),
            .in2(_gnd_net_),
            .in3(N__38138),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__49048),
            .ce(N__39574),
            .sr(N__48585));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_19_0  (
            .in0(N__39509),
            .in1(N__40440),
            .in2(_gnd_net_),
            .in3(N__38189),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__49041),
            .ce(N__39570),
            .sr(N__48593));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_19_1  (
            .in0(N__39536),
            .in1(N__40407),
            .in2(_gnd_net_),
            .in3(N__38186),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__49041),
            .ce(N__39570),
            .sr(N__48593));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_19_2  (
            .in0(N__39510),
            .in1(N__40377),
            .in2(_gnd_net_),
            .in3(N__38183),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__49041),
            .ce(N__39570),
            .sr(N__48593));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_19_3  (
            .in0(N__39537),
            .in1(N__40827),
            .in2(_gnd_net_),
            .in3(N__38180),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__49041),
            .ce(N__39570),
            .sr(N__48593));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_19_4  (
            .in0(N__39511),
            .in1(N__40803),
            .in2(_gnd_net_),
            .in3(N__38177),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__49041),
            .ce(N__39570),
            .sr(N__48593));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_19_5  (
            .in0(N__39538),
            .in1(N__40777),
            .in2(_gnd_net_),
            .in3(N__38174),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__49041),
            .ce(N__39570),
            .sr(N__48593));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_19_6  (
            .in0(N__39512),
            .in1(N__40747),
            .in2(_gnd_net_),
            .in3(N__38171),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__49041),
            .ce(N__39570),
            .sr(N__48593));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_19_7  (
            .in0(N__39539),
            .in1(N__40717),
            .in2(_gnd_net_),
            .in3(N__38168),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__49041),
            .ce(N__39570),
            .sr(N__48593));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_20_0  (
            .in0(N__39513),
            .in1(N__40692),
            .in2(_gnd_net_),
            .in3(N__38165),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__49033),
            .ce(N__39575),
            .sr(N__48603));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_20_1  (
            .in0(N__39534),
            .in1(N__40662),
            .in2(_gnd_net_),
            .in3(N__38288),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__49033),
            .ce(N__39575),
            .sr(N__48603));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_20_2  (
            .in0(N__39514),
            .in1(N__40620),
            .in2(_gnd_net_),
            .in3(N__38285),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__49033),
            .ce(N__39575),
            .sr(N__48603));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_20_3  (
            .in0(N__39535),
            .in1(N__41121),
            .in2(_gnd_net_),
            .in3(N__38282),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__49033),
            .ce(N__39575),
            .sr(N__48603));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_20_4  (
            .in0(N__39515),
            .in1(N__40639),
            .in2(_gnd_net_),
            .in3(N__38279),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__49033),
            .ce(N__39575),
            .sr(N__48603));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_20_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_20_5  (
            .in0(N__41140),
            .in1(N__39516),
            .in2(_gnd_net_),
            .in3(N__38276),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49033),
            .ce(N__39575),
            .sr(N__48603));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_21_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_21_0  (
            .in0(N__38259),
            .in1(N__38242),
            .in2(N__38201),
            .in3(N__38210),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_15_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_15_21_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_15_21_1  (
            .in0(N__38209),
            .in1(N__38260),
            .in2(N__38246),
            .in3(N__38197),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_15_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_15_21_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_15_21_2  (
            .in0(N__49742),
            .in1(N__49769),
            .in2(_gnd_net_),
            .in3(N__49576),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49028),
            .ce(N__48720),
            .sr(N__48612));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_15_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_15_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_15_21_3  (
            .in0(N__49574),
            .in1(N__48172),
            .in2(_gnd_net_),
            .in3(N__47006),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49028),
            .ce(N__48720),
            .sr(N__48612));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_15_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_15_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_15_21_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_15_21_7  (
            .in0(N__49575),
            .in1(N__47250),
            .in2(_gnd_net_),
            .in3(N__47227),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49028),
            .ce(N__48720),
            .sr(N__48612));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_22_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_22_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_22_0  (
            .in0(N__39710),
            .in1(N__47756),
            .in2(N__39771),
            .in3(N__47225),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_15_22_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_15_22_1 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_15_22_1  (
            .in0(N__50258),
            .in1(_gnd_net_),
            .in2(N__38312),
            .in3(N__43583),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_22_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_22_2  (
            .in0(N__39799),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49024),
            .ce(N__41094),
            .sr(N__48621));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_22_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_22_3  (
            .in0(N__39740),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49024),
            .ce(N__41094),
            .sr(N__48621));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_15_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_15_22_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_15_22_4  (
            .in0(N__47254),
            .in1(N__47226),
            .in2(_gnd_net_),
            .in3(N__49424),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_22_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_22_5  (
            .in0(N__47757),
            .in1(N__49425),
            .in2(_gnd_net_),
            .in3(N__47190),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_22_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_22_6  (
            .in0(N__39764),
            .in1(N__39330),
            .in2(_gnd_net_),
            .in3(N__49423),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_22_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_22_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_22_7  (
            .in0(N__49422),
            .in1(N__39303),
            .in2(_gnd_net_),
            .in3(N__39711),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_15_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_15_23_0 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_15_23_0  (
            .in0(N__38300),
            .in1(N__38472),
            .in2(N__38456),
            .in3(N__38342),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_15_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_15_23_3 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_15_23_3  (
            .in0(N__40864),
            .in1(N__40930),
            .in2(N__38390),
            .in3(N__38403),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_23_4 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_23_4  (
            .in0(N__38404),
            .in1(N__40865),
            .in2(N__40931),
            .in3(N__38388),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_23_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_23_5  (
            .in0(N__43558),
            .in1(N__43584),
            .in2(_gnd_net_),
            .in3(N__49534),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_15_24_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_15_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_15_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_15_24_0  (
            .in0(N__47090),
            .in1(N__47041),
            .in2(_gnd_net_),
            .in3(N__49628),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49015),
            .ce(N__48715),
            .sr(N__48634));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_15_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_15_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_15_24_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_15_24_2  (
            .in0(N__47501),
            .in1(N__48149),
            .in2(_gnd_net_),
            .in3(N__49625),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49015),
            .ce(N__48715),
            .sr(N__48634));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_15_24_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_15_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_15_24_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_15_24_3  (
            .in0(N__49624),
            .in1(N__39334),
            .in2(_gnd_net_),
            .in3(N__39773),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49015),
            .ce(N__48715),
            .sr(N__48634));
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_15_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_15_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_15_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_27_LC_15_24_4  (
            .in0(N__50260),
            .in1(N__50236),
            .in2(_gnd_net_),
            .in3(N__49626),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49015),
            .ce(N__48715),
            .sr(N__48634));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_15_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_15_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_15_24_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_15_24_6  (
            .in0(N__39307),
            .in1(N__39716),
            .in2(_gnd_net_),
            .in3(N__49627),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49015),
            .ce(N__48715),
            .sr(N__48634));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_25_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_25_0 .LUT_INIT=16'b0010101100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_25_0  (
            .in0(N__38627),
            .in1(N__38650),
            .in2(N__38675),
            .in3(N__41036),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_25_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_25_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_25_1  (
            .in0(N__41035),
            .in1(N__38674),
            .in2(N__38651),
            .in3(N__38626),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_15_25_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_15_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_15_25_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_15_25_4  (
            .in0(N__47191),
            .in1(N__47764),
            .in2(_gnd_net_),
            .in3(N__49577),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49013),
            .ce(N__48713),
            .sr(N__48638));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_26_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_26_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_26_6 .LUT_INIT=16'b1111010101110001;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_26_6  (
            .in0(N__40961),
            .in1(N__38557),
            .in2(N__38599),
            .in3(N__40888),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_15_27_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_15_27_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_15_27_2 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_15_27_2  (
            .in0(N__40887),
            .in1(N__38592),
            .in2(N__38558),
            .in3(N__40960),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_16_5_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_16_5_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_16_5_0 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_16_5_0  (
            .in0(N__39396),
            .in1(N__39610),
            .in2(_gnd_net_),
            .in3(N__39379),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49140),
            .ce(),
            .sr(N__48516));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_6_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_6_0  (
            .in0(N__44620),
            .in1(N__42451),
            .in2(N__44156),
            .in3(N__41516),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_16_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_16_6_1 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_16_6_1  (
            .in0(N__41167),
            .in1(N__44624),
            .in2(N__42473),
            .in3(N__46183),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_16_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_16_6_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_16_6_2  (
            .in0(N__44623),
            .in1(N__42447),
            .in2(N__45169),
            .in3(N__41572),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_6_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_6_4  (
            .in0(N__41863),
            .in1(N__46716),
            .in2(_gnd_net_),
            .in3(N__38973),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_16_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_16_6_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_16_6_6  (
            .in0(N__44621),
            .in1(N__42445),
            .in2(N__45323),
            .in3(N__38876),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_16_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_16_6_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_16_6_7  (
            .in0(N__42446),
            .in1(N__44622),
            .in2(N__45248),
            .in3(N__41495),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44222),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_7_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_7_1  (
            .in0(N__42459),
            .in1(N__44707),
            .in2(N__45827),
            .in3(N__41732),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45620),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_7_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_7_3  (
            .in0(N__41467),
            .in1(N__44708),
            .in2(N__42474),
            .in3(N__46861),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_16_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_16_7_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_16_7_4  (
            .in0(N__44705),
            .in1(N__42460),
            .in2(N__46112),
            .in3(N__42571),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_7_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_7_5  (
            .in0(N__42461),
            .in1(N__44706),
            .in2(N__45971),
            .in3(N__41653),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_7_7 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_7_7  (
            .in0(N__41627),
            .in1(N__44709),
            .in2(N__42475),
            .in3(N__46795),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__38834),
            .in2(N__38827),
            .in3(N__38828),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__41474),
            .in2(_gnd_net_),
            .in3(N__38804),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__41444),
            .in2(_gnd_net_),
            .in3(N__38801),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(N__38798),
            .in2(_gnd_net_),
            .in3(N__38792),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__41711),
            .in2(_gnd_net_),
            .in3(N__38789),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__41438),
            .in2(_gnd_net_),
            .in3(N__38786),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__38783),
            .in2(_gnd_net_),
            .in3(N__38777),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__41549),
            .in2(_gnd_net_),
            .in3(N__38774),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__38924),
            .in2(_gnd_net_),
            .in3(N__38882),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42662),
            .in3(N__38879),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42632),
            .in3(N__38855),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__42620),
            .in2(_gnd_net_),
            .in3(N__38852),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__41633),
            .in2(_gnd_net_),
            .in3(N__38849),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__42650),
            .in2(_gnd_net_),
            .in3(N__38846),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__42596),
            .in2(_gnd_net_),
            .in3(N__38843),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__39620),
            .in2(_gnd_net_),
            .in3(N__38840),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__39023),
            .in2(_gnd_net_),
            .in3(N__38837),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__42671),
            .in2(_gnd_net_),
            .in3(N__39005),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__42641),
            .in2(_gnd_net_),
            .in3(N__39002),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__42800),
            .in2(_gnd_net_),
            .in3(N__38999),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_10_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42791),
            .in3(N__38996),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__42818),
            .in2(_gnd_net_),
            .in3(N__38993),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_10_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42608),
            .in3(N__38990),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(N__42779),
            .in2(_gnd_net_),
            .in3(N__38954),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__42767),
            .in2(_gnd_net_),
            .in3(N__38951),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_11_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39014),
            .in3(N__38927),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__42809),
            .in2(_gnd_net_),
            .in3(N__39116),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__39029),
            .in2(_gnd_net_),
            .in3(N__39113),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__42584),
            .in2(_gnd_net_),
            .in3(N__39086),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39083),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_11_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_11_6  (
            .in0(N__42420),
            .in1(N__44759),
            .in2(N__46796),
            .in3(N__41623),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_16_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_16_11_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_16_11_7  (
            .in0(N__44758),
            .in1(N__42421),
            .in2(N__45896),
            .in3(N__42547),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46406),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46028),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46562),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46094),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_13_1 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_13_1  (
            .in0(N__39380),
            .in1(N__39407),
            .in2(_gnd_net_),
            .in3(N__39611),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_202_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39405),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_14_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_14_2  (
            .in0(N__39406),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39375),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_201_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_16_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_16_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_16_15_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_16_15_4  (
            .in0(N__39338),
            .in1(N__39772),
            .in2(_gnd_net_),
            .in3(N__49582),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49075),
            .ce(N__49952),
            .sr(N__48548));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_16_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_16_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_16_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_16_15_6  (
            .in0(N__39715),
            .in1(N__39308),
            .in2(_gnd_net_),
            .in3(N__49583),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49075),
            .ce(N__49952),
            .sr(N__48548));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_16_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_16_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_16_15_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_16_15_7  (
            .in0(N__49581),
            .in1(N__39281),
            .in2(_gnd_net_),
            .in3(N__40277),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49075),
            .ce(N__49952),
            .sr(N__48548));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_16_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_16_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_16_16_0 .LUT_INIT=16'b1111001101000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_16_16_0  (
            .in0(N__43103),
            .in1(N__39670),
            .in2(N__50108),
            .in3(N__39251),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49068),
            .ce(),
            .sr(N__48556));
    defparam \phase_controller_inst1.T01_LC_16_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_16_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_16_16_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst1.T01_LC_16_16_6  (
            .in0(N__39127),
            .in1(N__39227),
            .in2(_gnd_net_),
            .in3(N__39173),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49068),
            .ce(),
            .sr(N__48556));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_16_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_16_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_16_16_7 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_16_16_7  (
            .in0(N__39669),
            .in1(N__39878),
            .in2(N__43091),
            .in3(N__50052),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49068),
            .ce(),
            .sr(N__48556));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_17_2 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_17_2  (
            .in0(N__39679),
            .in1(N__50134),
            .in2(_gnd_net_),
            .in3(N__50098),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_17_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39683),
            .in3(N__39873),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_LC_16_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_16_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_16_17_4 .LUT_INIT=16'b1000101011111010;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_16_17_4  (
            .in0(N__39680),
            .in1(N__43102),
            .in2(N__39671),
            .in3(N__50099),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49062),
            .ce(),
            .sr(N__48567));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_16_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_16_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__39665),
            .in2(_gnd_net_),
            .in3(N__39874),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_18_3 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_18_3  (
            .in0(N__39635),
            .in1(N__39650),
            .in2(N__43703),
            .in3(N__43734),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_16_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_16_18_4 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_16_18_4  (
            .in0(N__39649),
            .in1(N__39633),
            .in2(N__43735),
            .in3(N__43698),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_16_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_16_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_16_18_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_30_LC_16_18_5  (
            .in0(N__40915),
            .in1(N__43873),
            .in2(N__49623),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49056),
            .ce(N__49994),
            .sr(N__48578));
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_16_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_16_18_6 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_16_18_6  (
            .in0(N__39648),
            .in1(N__39634),
            .in2(N__43736),
            .in3(N__43699),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_16_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_16_18_7 .LUT_INIT=16'b1111110101011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_16_18_7  (
            .in0(N__50101),
            .in1(N__43126),
            .in2(N__39623),
            .in3(N__43115),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_19_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_19_0  (
            .in0(N__39839),
            .in1(N__39809),
            .in2(N__43463),
            .in3(N__43440),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_19_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_19_1  (
            .in0(N__39808),
            .in1(N__43461),
            .in2(N__43442),
            .in3(N__39838),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_19_2  (
            .in0(N__43524),
            .in1(N__39856),
            .in2(_gnd_net_),
            .in3(N__49530),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(elapsed_time_ns_1_RNI14DN9_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_16_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_16_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_16_19_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_23_LC_16_19_3  (
            .in0(N__49533),
            .in1(_gnd_net_),
            .in2(N__39842),
            .in3(N__43525),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49049),
            .ce(N__50006),
            .sr(N__48586));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_19_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_19_4  (
            .in0(N__43497),
            .in1(N__39823),
            .in2(_gnd_net_),
            .in3(N__49531),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(elapsed_time_ns_1_RNI03DN9_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_16_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_16_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_16_19_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_22_LC_16_19_5  (
            .in0(N__49532),
            .in1(_gnd_net_),
            .in2(N__39812),
            .in3(N__43498),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49049),
            .ce(N__50006),
            .sr(N__48586));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_20_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__40354),
            .in2(N__39800),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49042),
            .ce(N__41087),
            .sr(N__48594));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(N__39739),
            .in2(N__40333),
            .in3(N__39686),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49042),
            .ce(N__41087),
            .sr(N__48594));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__40355),
            .in2(N__40304),
            .in3(N__40337),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49042),
            .ce(N__41087),
            .sr(N__48594));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(N__40231),
            .in2(N__40334),
            .in3(N__40307),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49042),
            .ce(N__41087),
            .sr(N__48594));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__40303),
            .in2(N__40168),
            .in3(N__40235),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49042),
            .ce(N__41087),
            .sr(N__48594));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(N__40232),
            .in2(N__40099),
            .in3(N__40172),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49042),
            .ce(N__41087),
            .sr(N__48594));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__40024),
            .in2(N__40169),
            .in3(N__40103),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49042),
            .ce(N__41087),
            .sr(N__48594));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(N__39952),
            .in2(N__40100),
            .in3(N__40034),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49042),
            .ce(N__41087),
            .sr(N__48594));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__40597),
            .in2(N__40031),
            .in3(N__39962),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49034),
            .ce(N__41083),
            .sr(N__48604));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__40576),
            .in2(N__39959),
            .in3(N__39881),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49034),
            .ce(N__41083),
            .sr(N__48604));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__40598),
            .in2(N__40556),
            .in3(N__40580),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49034),
            .ce(N__41083),
            .sr(N__48604));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__40577),
            .in2(N__40529),
            .in3(N__40559),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49034),
            .ce(N__41083),
            .sr(N__48604));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__40555),
            .in2(N__40501),
            .in3(N__40532),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49034),
            .ce(N__41083),
            .sr(N__48604));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(N__40528),
            .in2(N__40474),
            .in3(N__40505),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49034),
            .ce(N__41083),
            .sr(N__48604));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(N__40441),
            .in2(N__40502),
            .in3(N__40478),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49034),
            .ce(N__41083),
            .sr(N__48604));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(N__40414),
            .in2(N__40475),
            .in3(N__40451),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49034),
            .ce(N__41083),
            .sr(N__48604));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__40378),
            .in2(N__40448),
            .in3(N__40421),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49029),
            .ce(N__41095),
            .sr(N__48613));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(N__40828),
            .in2(N__40418),
            .in3(N__40385),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49029),
            .ce(N__41095),
            .sr(N__48613));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(N__40804),
            .in2(N__40382),
            .in3(N__40358),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49029),
            .ce(N__41095),
            .sr(N__48613));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__40783),
            .in2(N__40832),
            .in3(N__40808),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49029),
            .ce(N__41095),
            .sr(N__48613));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(N__40805),
            .in2(N__40759),
            .in3(N__40787),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49029),
            .ce(N__41095),
            .sr(N__48613));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(N__40784),
            .in2(N__40729),
            .in3(N__40763),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49029),
            .ce(N__41095),
            .sr(N__48613));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_22_6  (
            .in0(_gnd_net_),
            .in1(N__40693),
            .in2(N__40760),
            .in3(N__40733),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49029),
            .ce(N__41095),
            .sr(N__48613));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_22_7  (
            .in0(_gnd_net_),
            .in1(N__40663),
            .in2(N__40730),
            .in3(N__40703),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49029),
            .ce(N__41095),
            .sr(N__48613));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(N__40621),
            .in2(N__40700),
            .in3(N__40673),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49025),
            .ce(N__41096),
            .sr(N__48622));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_23_1  (
            .in0(_gnd_net_),
            .in1(N__41122),
            .in2(N__40670),
            .in3(N__40643),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49025),
            .ce(N__41096),
            .sr(N__48622));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(N__40640),
            .in2(N__40625),
            .in3(N__40601),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49025),
            .ce(N__41096),
            .sr(N__48622));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(N__41144),
            .in2(N__41126),
            .in3(N__41102),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49025),
            .ce(N__41096),
            .sr(N__48622));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41099),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49025),
            .ce(N__41096),
            .sr(N__48622));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_16_24_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_16_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_16_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_16_24_0  (
            .in0(N__48072),
            .in1(N__48221),
            .in2(_gnd_net_),
            .in3(N__49568),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49020),
            .ce(N__48718),
            .sr(N__48628));
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_16_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_16_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_16_24_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_31_LC_16_24_1  (
            .in0(N__49567),
            .in1(N__41007),
            .in2(_gnd_net_),
            .in3(N__40991),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49020),
            .ce(N__48718),
            .sr(N__48628));
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_16_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_16_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_16_24_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_29_LC_16_24_2  (
            .in0(N__43616),
            .in1(N__43895),
            .in2(_gnd_net_),
            .in3(N__49570),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49020),
            .ce(N__48718),
            .sr(N__48628));
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_16_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_16_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_16_24_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_30_LC_16_24_4  (
            .in0(N__40919),
            .in1(N__43866),
            .in2(_gnd_net_),
            .in3(N__49571),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49020),
            .ce(N__48718),
            .sr(N__48628));
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_16_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_16_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_16_24_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_28_LC_16_24_6  (
            .in0(N__43585),
            .in1(N__43554),
            .in2(_gnd_net_),
            .in3(N__49569),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49020),
            .ce(N__48718),
            .sr(N__48628));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_16_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_16_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_16_25_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_16_25_5  (
            .in0(N__47631),
            .in1(N__47890),
            .in2(_gnd_net_),
            .in3(N__49554),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49016),
            .ce(N__48716),
            .sr(N__48635));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_17_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_17_7_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_17_7_0  (
            .in0(N__41425),
            .in1(N__44704),
            .in2(N__42476),
            .in3(N__45622),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_7_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_7_1  (
            .in0(N__45621),
            .in1(N__41855),
            .in2(_gnd_net_),
            .in3(N__41424),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_7_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_7_2  (
            .in0(N__41853),
            .in1(N__44298),
            .in2(_gnd_net_),
            .in3(N__41400),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_7_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_7_4  (
            .in0(N__41852),
            .in1(N__41379),
            .in2(_gnd_net_),
            .in3(N__41363),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_7_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_7_5  (
            .in0(N__45687),
            .in1(N__41854),
            .in2(_gnd_net_),
            .in3(N__41325),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_7_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_7_6  (
            .in0(N__41856),
            .in1(N__45549),
            .in2(_gnd_net_),
            .in3(N__41301),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_17_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_17_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41285),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_8_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_8_1  (
            .in0(N__46245),
            .in1(N__41861),
            .in2(_gnd_net_),
            .in3(N__41199),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_8_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_8_2  (
            .in0(N__41857),
            .in1(N__41181),
            .in2(_gnd_net_),
            .in3(N__44356),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_8_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_8_3  (
            .in0(N__46176),
            .in1(N__41862),
            .in2(_gnd_net_),
            .in3(N__41160),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_8_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_8_4  (
            .in0(N__41860),
            .in1(N__45151),
            .in2(_gnd_net_),
            .in3(N__41565),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45548),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_8_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_8_6  (
            .in0(N__41858),
            .in1(_gnd_net_),
            .in2(N__44223),
            .in3(N__41532),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_8_7 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_8_7  (
            .in0(N__41508),
            .in1(N__41859),
            .in2(_gnd_net_),
            .in3(N__44137),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_9_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_9_0  (
            .in0(N__45231),
            .in1(N__41844),
            .in2(_gnd_net_),
            .in3(N__41490),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_9_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__44355),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_9_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_9_2  (
            .in0(N__46854),
            .in1(N__41846),
            .in2(_gnd_net_),
            .in3(N__41460),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44288),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_9_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_9_4  (
            .in0(N__45677),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_9_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_9_5  (
            .in0(N__41843),
            .in1(N__45393),
            .in2(_gnd_net_),
            .in3(N__41748),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_9_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_9_6  (
            .in0(N__45819),
            .in1(N__41845),
            .in2(_gnd_net_),
            .in3(N__41727),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44136),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_10_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_10_0  (
            .in0(N__44725),
            .in1(N__46641),
            .in2(_gnd_net_),
            .in3(N__41694),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_10_1 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_10_1  (
            .in0(N__41803),
            .in1(N__41676),
            .in2(_gnd_net_),
            .in3(N__46035),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_10_2 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_10_2  (
            .in0(N__45963),
            .in1(N__41646),
            .in2(_gnd_net_),
            .in3(N__41804),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_10_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_10_3  (
            .in0(N__45144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_10_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_10_4  (
            .in0(N__46782),
            .in1(N__41806),
            .in2(_gnd_net_),
            .in3(N__41622),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_10_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_10_5  (
            .in0(N__46497),
            .in1(N__44726),
            .in2(_gnd_net_),
            .in3(N__41598),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_10_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_10_6  (
            .in0(N__46101),
            .in1(N__41802),
            .in2(_gnd_net_),
            .in3(N__42570),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_10_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_10_7  (
            .in0(N__41805),
            .in1(_gnd_net_),
            .in2(N__45891),
            .in3(N__42546),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_11_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_11_1  (
            .in0(N__46408),
            .in1(N__44756),
            .in2(N__42515),
            .in3(N__42399),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_11_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_11_2  (
            .in0(N__44753),
            .in1(N__46407),
            .in2(_gnd_net_),
            .in3(N__42510),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_11_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__44757),
            .in2(_gnd_net_),
            .in3(N__42398),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_11_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_11_4  (
            .in0(N__44754),
            .in1(N__45748),
            .in2(N__42465),
            .in3(N__41878),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_11_5 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_11_5  (
            .in0(N__45749),
            .in1(N__44755),
            .in2(N__41879),
            .in3(N__42403),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_11_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_11_6  (
            .in0(N__41807),
            .in1(N__45747),
            .in2(_gnd_net_),
            .in3(N__41874),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47121),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49117),
            .ce(N__47164),
            .sr(N__48523));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45945),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45375),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46228),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45873),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_17_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_17_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45294),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45221),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46772),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46158),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46302),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46836),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46478),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45800),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45739),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46697),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46623),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_17_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_17_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42758),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__47207),
            .in2(N__42689),
            .in3(N__43083),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__47738),
            .in2(N__42680),
            .in3(N__43058),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__42947),
            .in2(N__42941),
            .in3(N__43033),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__42932),
            .in2(N__42926),
            .in3(N__43313),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__42917),
            .in2(N__47336),
            .in3(N__43295),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_15_5  (
            .in0(N__43277),
            .in1(N__47018),
            .in2(N__42911),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__42902),
            .in2(N__42896),
            .in3(N__43259),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__42884),
            .in2(N__42872),
            .in3(N__43241),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__42860),
            .in2(N__42848),
            .in3(N__43223),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__42839),
            .in2(N__42827),
            .in3(N__43205),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__43013),
            .in2(N__43001),
            .in3(N__43184),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__42992),
            .in2(N__42980),
            .in3(N__43403),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__43820),
            .in2(N__42971),
            .in3(N__43385),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_16_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_16_5  (
            .in0(N__43367),
            .in1(N__46892),
            .in2(N__42962),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__42953),
            .in2(N__47615),
            .in3(N__43349),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__47012),
            .in2(N__46925),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__47510),
            .in2(N__47558),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__47318),
            .in2(N__47270),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__43166),
            .in2(N__43154),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__47402),
            .in2(N__47462),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__48191),
            .in2(N__47975),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__43625),
            .in2(N__43676),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__43139),
            .in2(N__43133),
            .in3(N__43109),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43106),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__43090),
            .in2(N__43067),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_17_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_17_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_17_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_17_18_1  (
            .in0(N__49998),
            .in1(N__43057),
            .in2(_gnd_net_),
            .in3(N__43043),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49063),
            .ce(),
            .sr(N__48568));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_17_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_17_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_17_18_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_17_18_2  (
            .in0(N__49975),
            .in1(N__43040),
            .in2(N__43034),
            .in3(N__43016),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49063),
            .ce(),
            .sr(N__48568));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_17_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_17_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_17_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_17_18_3  (
            .in0(N__49999),
            .in1(N__43312),
            .in2(_gnd_net_),
            .in3(N__43298),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49063),
            .ce(),
            .sr(N__48568));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_17_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_17_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_17_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_17_18_4  (
            .in0(N__49976),
            .in1(N__43294),
            .in2(_gnd_net_),
            .in3(N__43280),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49063),
            .ce(),
            .sr(N__48568));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_17_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_17_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_17_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_17_18_5  (
            .in0(N__50000),
            .in1(N__43276),
            .in2(_gnd_net_),
            .in3(N__43262),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49063),
            .ce(),
            .sr(N__48568));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_17_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_17_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_17_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_17_18_6  (
            .in0(N__49977),
            .in1(N__43258),
            .in2(_gnd_net_),
            .in3(N__43244),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49063),
            .ce(),
            .sr(N__48568));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_17_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_17_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_17_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_17_18_7  (
            .in0(N__50001),
            .in1(N__43240),
            .in2(_gnd_net_),
            .in3(N__43226),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49063),
            .ce(),
            .sr(N__48568));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_17_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_17_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_17_19_0  (
            .in0(N__49981),
            .in1(N__43222),
            .in2(_gnd_net_),
            .in3(N__43208),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49057),
            .ce(),
            .sr(N__48579));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_17_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_17_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_17_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_17_19_1  (
            .in0(N__49961),
            .in1(N__43201),
            .in2(_gnd_net_),
            .in3(N__43187),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49057),
            .ce(),
            .sr(N__48579));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_17_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_17_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_17_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_17_19_2  (
            .in0(N__49978),
            .in1(N__43183),
            .in2(_gnd_net_),
            .in3(N__43169),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49057),
            .ce(),
            .sr(N__48579));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_17_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_17_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_17_19_3  (
            .in0(N__49962),
            .in1(N__43402),
            .in2(_gnd_net_),
            .in3(N__43388),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49057),
            .ce(),
            .sr(N__48579));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_17_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_17_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_17_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_17_19_4  (
            .in0(N__49979),
            .in1(N__43384),
            .in2(_gnd_net_),
            .in3(N__43370),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49057),
            .ce(),
            .sr(N__48579));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_17_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_17_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_17_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_17_19_5  (
            .in0(N__49963),
            .in1(N__43366),
            .in2(_gnd_net_),
            .in3(N__43352),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49057),
            .ce(),
            .sr(N__48579));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_17_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_17_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_17_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_17_19_6  (
            .in0(N__49980),
            .in1(N__43345),
            .in2(_gnd_net_),
            .in3(N__43331),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49057),
            .ce(),
            .sr(N__48579));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_17_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_17_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_17_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_17_19_7  (
            .in0(N__49964),
            .in1(N__46948),
            .in2(_gnd_net_),
            .in3(N__43328),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49057),
            .ce(),
            .sr(N__48579));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_17_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_17_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_17_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_17_20_0  (
            .in0(N__49953),
            .in1(N__46975),
            .in2(_gnd_net_),
            .in3(N__43325),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49050),
            .ce(),
            .sr(N__48587));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_17_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_17_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_17_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_17_20_1  (
            .in0(N__50048),
            .in1(N__47543),
            .in2(_gnd_net_),
            .in3(N__43322),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49050),
            .ce(),
            .sr(N__48587));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_17_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_17_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_17_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_17_20_2  (
            .in0(N__49954),
            .in1(N__47527),
            .in2(_gnd_net_),
            .in3(N__43319),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49050),
            .ce(),
            .sr(N__48587));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_17_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_17_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_17_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_17_20_3  (
            .in0(N__50049),
            .in1(N__47310),
            .in2(_gnd_net_),
            .in3(N__43316),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49050),
            .ce(),
            .sr(N__48587));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_17_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_17_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_17_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_17_20_4  (
            .in0(N__49955),
            .in1(N__47286),
            .in2(_gnd_net_),
            .in3(N__43466),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49050),
            .ce(),
            .sr(N__48587));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_17_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_17_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_17_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_17_20_5  (
            .in0(N__50050),
            .in1(N__43462),
            .in2(_gnd_net_),
            .in3(N__43445),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49050),
            .ce(),
            .sr(N__48587));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_17_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_17_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_17_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_17_20_6  (
            .in0(N__49956),
            .in1(N__43441),
            .in2(_gnd_net_),
            .in3(N__43424),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49050),
            .ce(),
            .sr(N__48587));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_17_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_17_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_17_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_17_20_7  (
            .in0(N__50051),
            .in1(N__47418),
            .in2(_gnd_net_),
            .in3(N__43421),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49050),
            .ce(),
            .sr(N__48587));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_17_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_17_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_17_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_17_21_0  (
            .in0(N__49957),
            .in1(N__47445),
            .in2(_gnd_net_),
            .in3(N__43418),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49043),
            .ce(),
            .sr(N__48595));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_17_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_17_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_17_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_17_21_1  (
            .in0(N__50053),
            .in1(N__48005),
            .in2(_gnd_net_),
            .in3(N__43415),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49043),
            .ce(),
            .sr(N__48595));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_17_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_17_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_17_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_17_21_2  (
            .in0(N__49958),
            .in1(N__47990),
            .in2(_gnd_net_),
            .in3(N__43412),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49043),
            .ce(),
            .sr(N__48595));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_17_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_17_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_17_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_17_21_3  (
            .in0(N__50054),
            .in1(N__43661),
            .in2(_gnd_net_),
            .in3(N__43409),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49043),
            .ce(),
            .sr(N__48595));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_17_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_17_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_17_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_17_21_4  (
            .in0(N__49959),
            .in1(N__43641),
            .in2(_gnd_net_),
            .in3(N__43406),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49043),
            .ce(),
            .sr(N__48595));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_17_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_17_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_17_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_17_21_5  (
            .in0(N__50055),
            .in1(N__43727),
            .in2(_gnd_net_),
            .in3(N__43709),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49043),
            .ce(),
            .sr(N__48595));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_17_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_17_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_17_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_17_21_6  (
            .in0(N__49960),
            .in1(N__43690),
            .in2(_gnd_net_),
            .in3(N__43706),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49043),
            .ce(),
            .sr(N__48595));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_17_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_17_22_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_17_22_0  (
            .in0(N__43659),
            .in1(N__43642),
            .in2(N__43598),
            .in3(N__43538),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_17_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_17_22_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_17_22_1  (
            .in0(N__43537),
            .in1(N__43660),
            .in2(N__43646),
            .in3(N__43594),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_17_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_17_22_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_17_22_2  (
            .in0(N__43893),
            .in1(N__43612),
            .in2(_gnd_net_),
            .in3(N__49454),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_17_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_17_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_17_22_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_29_LC_17_22_3  (
            .in0(N__49456),
            .in1(_gnd_net_),
            .in2(N__43601),
            .in3(N__43894),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49035),
            .ce(N__50032),
            .sr(N__48605));
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_17_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_17_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_17_22_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_28_LC_17_22_7  (
            .in0(N__49455),
            .in1(N__43586),
            .in2(_gnd_net_),
            .in3(N__43562),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49035),
            .ce(N__50032),
            .sr(N__48605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_23_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_23_3  (
            .in0(N__43515),
            .in1(N__43482),
            .in2(N__47678),
            .in3(N__47356),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_23_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_23_4  (
            .in0(N__43892),
            .in1(N__50162),
            .in2(N__47948),
            .in3(N__43862),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_17_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_17_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_17_23_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_17_23_6  (
            .in0(N__43841),
            .in1(N__49616),
            .in2(_gnd_net_),
            .in3(N__47808),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49030),
            .ce(N__50033),
            .sr(N__48614));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_17_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_17_24_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_17_24_0  (
            .in0(N__49637),
            .in1(N__48143),
            .in2(_gnd_net_),
            .in3(N__47493),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_24_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_24_1  (
            .in0(N__47635),
            .in1(N__47886),
            .in2(_gnd_net_),
            .in3(N__49636),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_17_24_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_17_24_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_17_24_4  (
            .in0(N__49638),
            .in1(N__50259),
            .in2(_gnd_net_),
            .in3(N__50235),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_24_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_24_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_24_6  (
            .in0(N__49635),
            .in1(N__47094),
            .in2(_gnd_net_),
            .in3(N__47040),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_18_7_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_18_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_18_7_0  (
            .in0(_gnd_net_),
            .in1(N__43808),
            .in2(N__43772),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_7_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_18_7_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_18_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_18_7_1  (
            .in0(_gnd_net_),
            .in1(N__45075),
            .in2(N__43751),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_18_7_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_18_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_18_7_2  (
            .in0(_gnd_net_),
            .in1(N__43742),
            .in2(N__45096),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_18_7_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_18_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_18_7_3  (
            .in0(_gnd_net_),
            .in1(N__45079),
            .in2(N__43976),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_18_7_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_18_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_18_7_4  (
            .in0(_gnd_net_),
            .in1(N__43967),
            .in2(N__45097),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_18_7_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_18_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_18_7_5  (
            .in0(_gnd_net_),
            .in1(N__45083),
            .in2(N__43961),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_18_7_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_18_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_18_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_18_7_6  (
            .in0(_gnd_net_),
            .in1(N__43952),
            .in2(N__45098),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_18_7_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_18_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_18_7_7  (
            .in0(_gnd_net_),
            .in1(N__45087),
            .in2(N__43946),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_18_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_18_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_18_8_0  (
            .in0(_gnd_net_),
            .in1(N__44965),
            .in2(N__43937),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_8_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_18_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_18_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_18_8_1  (
            .in0(_gnd_net_),
            .in1(N__43928),
            .in2(N__45039),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_18_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_18_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_18_8_2  (
            .in0(_gnd_net_),
            .in1(N__44953),
            .in2(N__43913),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_18_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_18_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(N__43904),
            .in2(N__45036),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_18_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_18_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(N__44957),
            .in2(N__44036),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_18_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_18_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(N__44027),
            .in2(N__45037),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_18_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_18_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_18_8_6  (
            .in0(_gnd_net_),
            .in1(N__44961),
            .in2(N__44021),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_18_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_18_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_18_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_18_8_7  (
            .in0(_gnd_net_),
            .in1(N__44012),
            .in2(N__45038),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_18_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_18_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_18_9_0  (
            .in0(_gnd_net_),
            .in1(N__45059),
            .in2(N__44006),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_9_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_18_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_18_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_18_9_1  (
            .in0(_gnd_net_),
            .in1(N__43997),
            .in2(N__45092),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_18_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_18_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_18_9_2  (
            .in0(_gnd_net_),
            .in1(N__45063),
            .in2(N__43991),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_18_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_18_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_18_9_3  (
            .in0(_gnd_net_),
            .in1(N__43982),
            .in2(N__45093),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_18_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_18_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_18_9_4  (
            .in0(_gnd_net_),
            .in1(N__45067),
            .in2(N__44111),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_18_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_18_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_18_9_5  (
            .in0(_gnd_net_),
            .in1(N__44102),
            .in2(N__45094),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_18_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_18_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_18_9_6  (
            .in0(_gnd_net_),
            .in1(N__45071),
            .in2(N__44093),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_18_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_18_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_18_9_7  (
            .in0(_gnd_net_),
            .in1(N__44084),
            .in2(N__45095),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_18_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_18_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__45046),
            .in2(N__44078),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_18_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_18_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(N__44063),
            .in2(N__45089),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_18_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_18_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_18_10_2  (
            .in0(_gnd_net_),
            .in1(N__45050),
            .in2(N__44057),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_18_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_18_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(N__44042),
            .in2(N__45090),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_18_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_18_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_18_10_4  (
            .in0(_gnd_net_),
            .in1(N__45054),
            .in2(N__45119),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_18_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_18_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(N__45107),
            .in2(N__45091),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_18_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_18_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_18_10_6  (
            .in0(_gnd_net_),
            .in1(N__45058),
            .in2(N__44774),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_10_7  (
            .in0(_gnd_net_),
            .in1(N__44727),
            .in2(_gnd_net_),
            .in3(N__44474),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__44392),
            .in2(N__44260),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49124),
            .ce(N__47167),
            .sr(N__48520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_11_1  (
            .in0(_gnd_net_),
            .in1(N__44336),
            .in2(N__44182),
            .in3(N__44264),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49124),
            .ce(N__47167),
            .sr(N__48520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__45721),
            .in2(N__44261),
            .in3(N__44186),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49124),
            .ce(N__47167),
            .sr(N__48520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(N__45646),
            .in2(N__44183),
            .in3(N__44114),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49124),
            .ce(N__47167),
            .sr(N__48520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__45583),
            .in2(N__45725),
            .in3(N__45650),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49124),
            .ce(N__47167),
            .sr(N__48520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__45647),
            .in2(N__45505),
            .in3(N__45587),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49124),
            .ce(N__47167),
            .sr(N__48520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__45584),
            .in2(N__45439),
            .in3(N__45509),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49124),
            .ce(N__47167),
            .sr(N__48520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(N__45352),
            .in2(N__45506),
            .in3(N__45443),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49124),
            .ce(N__47167),
            .sr(N__48520));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__45271),
            .in2(N__45440),
            .in3(N__45359),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49118),
            .ce(N__47165),
            .sr(N__48524));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__45193),
            .in2(N__45356),
            .in3(N__45278),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49118),
            .ce(N__47165),
            .sr(N__48524));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_12_2  (
            .in0(_gnd_net_),
            .in1(N__46279),
            .in2(N__45275),
            .in3(N__45200),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49118),
            .ce(N__47165),
            .sr(N__48524));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_12_3  (
            .in0(_gnd_net_),
            .in1(N__46213),
            .in2(N__45197),
            .in3(N__45122),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49118),
            .ce(N__47165),
            .sr(N__48524));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_12_4  (
            .in0(_gnd_net_),
            .in1(N__46135),
            .in2(N__46283),
            .in3(N__46217),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49118),
            .ce(N__47165),
            .sr(N__48524));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(N__46214),
            .in2(N__46063),
            .in3(N__46142),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49118),
            .ce(N__47165),
            .sr(N__48524));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(N__45994),
            .in2(N__46139),
            .in3(N__46067),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49118),
            .ce(N__47165),
            .sr(N__48524));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_12_7  (
            .in0(_gnd_net_),
            .in1(N__45919),
            .in2(N__46064),
            .in3(N__46004),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49118),
            .ce(N__47165),
            .sr(N__48524));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__45850),
            .in2(N__46001),
            .in3(N__45929),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49108),
            .ce(N__47162),
            .sr(N__48526));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__45772),
            .in2(N__45926),
            .in3(N__45857),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49108),
            .ce(N__47162),
            .sr(N__48526));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_13_2  (
            .in0(_gnd_net_),
            .in1(N__46885),
            .in2(N__45854),
            .in3(N__45779),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49108),
            .ce(N__47162),
            .sr(N__48526));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__46816),
            .in2(N__45776),
            .in3(N__45728),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49108),
            .ce(N__47162),
            .sr(N__48526));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__46886),
            .in2(N__46750),
            .in3(N__46820),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49108),
            .ce(N__47162),
            .sr(N__48526));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__46817),
            .in2(N__46672),
            .in3(N__46754),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49108),
            .ce(N__47162),
            .sr(N__48526));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(N__46597),
            .in2(N__46751),
            .in3(N__46676),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49108),
            .ce(N__47162),
            .sr(N__48526));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(N__46528),
            .in2(N__46673),
            .in3(N__46607),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49108),
            .ce(N__47162),
            .sr(N__48526));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__46432),
            .in2(N__46604),
            .in3(N__46538),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49101),
            .ce(N__47161),
            .sr(N__48530));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__46351),
            .in2(N__46535),
            .in3(N__46457),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49101),
            .ce(N__47161),
            .sr(N__48530));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__46454),
            .in2(N__46436),
            .in3(N__46376),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49101),
            .ce(N__47161),
            .sr(N__48530));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__46373),
            .in2(N__46355),
            .in3(N__46286),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49101),
            .ce(N__47161),
            .sr(N__48530));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47138),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_18_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_18_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_18_15_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_18_15_0  (
            .in0(N__47096),
            .in1(N__47048),
            .in2(_gnd_net_),
            .in3(N__49640),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49093),
            .ce(N__50066),
            .sr(N__48536));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_16_0 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_16_0  (
            .in0(N__46982),
            .in1(N__47570),
            .in2(N__46961),
            .in3(N__46934),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_16_2  (
            .in0(N__49584),
            .in1(N__48178),
            .in2(_gnd_net_),
            .in3(N__46996),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(elapsed_time_ns_1_RNI46CN9_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_18_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_18_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_18_16_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_18_16_3  (
            .in0(N__48179),
            .in1(_gnd_net_),
            .in2(N__46985),
            .in3(N__49587),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49084),
            .ce(N__50034),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_18_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_18_16_4 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_18_16_4  (
            .in0(N__46981),
            .in1(N__47569),
            .in2(N__46960),
            .in3(N__46933),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_18_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_18_16_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_18_16_5  (
            .in0(N__47851),
            .in1(N__49585),
            .in2(_gnd_net_),
            .in3(N__46906),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(elapsed_time_ns_1_RNI13CN9_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_18_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_18_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_18_16_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_18_16_6  (
            .in0(N__49586),
            .in1(_gnd_net_),
            .in2(N__46895),
            .in3(N__47852),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49084),
            .ce(N__50034),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_17_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_17_0  (
            .in0(N__47425),
            .in1(N__47453),
            .in2(N__47726),
            .in3(N__47345),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_18_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_18_17_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_18_17_1  (
            .in0(N__47344),
            .in1(N__47452),
            .in2(N__47429),
            .in3(N__47722),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_18_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_18_17_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_18_17_4  (
            .in0(N__47376),
            .in1(N__47392),
            .in2(_gnd_net_),
            .in3(N__49629),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(elapsed_time_ns_1_RNI25DN9_0_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_18_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_18_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_18_17_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_24_LC_18_17_5  (
            .in0(N__49630),
            .in1(_gnd_net_),
            .in2(N__47381),
            .in3(N__47377),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49076),
            .ce(N__50062),
            .sr(N__48549));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_18_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_18_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_18_17_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_18_17_6  (
            .in0(N__49714),
            .in1(N__49666),
            .in2(_gnd_net_),
            .in3(N__49631),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49076),
            .ce(N__50062),
            .sr(N__48549));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_18_0 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_18_0  (
            .in0(N__47579),
            .in1(N__47312),
            .in2(N__47294),
            .in3(N__47648),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_18_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_18_4  (
            .in0(N__47578),
            .in1(N__47311),
            .in2(N__47293),
            .in3(N__47647),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_18_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_18_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_18_18_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_18_18_6  (
            .in0(N__47258),
            .in1(N__47234),
            .in2(_gnd_net_),
            .in3(N__49619),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49069),
            .ce(N__49990),
            .sr(N__48557));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_18_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_18_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_18_18_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_18_18_7  (
            .in0(N__49618),
            .in1(N__47195),
            .in2(_gnd_net_),
            .in3(N__47768),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49069),
            .ce(N__49990),
            .sr(N__48557));
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_18_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_18_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_18_19_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_25_LC_18_19_1  (
            .in0(N__47914),
            .in1(N__47960),
            .in2(_gnd_net_),
            .in3(N__49592),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49064),
            .ce(N__50005),
            .sr(N__48569));
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_18_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_18_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_18_19_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_21_LC_18_19_3  (
            .in0(N__47711),
            .in1(N__47687),
            .in2(_gnd_net_),
            .in3(N__49591),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49064),
            .ce(N__50005),
            .sr(N__48569));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_18_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_18_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_18_19_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_18_19_5  (
            .in0(N__47639),
            .in1(N__47891),
            .in2(_gnd_net_),
            .in3(N__49589),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49064),
            .ce(N__50005),
            .sr(N__48569));
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_18_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_18_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_18_19_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_20_LC_18_19_6  (
            .in0(N__49588),
            .in1(N__47603),
            .in2(_gnd_net_),
            .in3(N__48111),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49064),
            .ce(N__50005),
            .sr(N__48569));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_18_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_18_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_18_19_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_18_19_7  (
            .in0(N__49741),
            .in1(N__49778),
            .in2(_gnd_net_),
            .in3(N__49590),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49064),
            .ce(N__50005),
            .sr(N__48569));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_20_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_20_0  (
            .in0(N__47541),
            .in1(N__47523),
            .in2(N__47474),
            .in3(N__48200),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_20_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_20_1  (
            .in0(N__48199),
            .in1(N__47542),
            .in2(N__47528),
            .in3(N__47470),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_18_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_18_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_18_20_3  (
            .in0(N__49615),
            .in1(N__47500),
            .in2(_gnd_net_),
            .in3(N__48148),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49058),
            .ce(N__50047),
            .sr(N__48580));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_20_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_20_6  (
            .in0(N__48073),
            .in1(N__48214),
            .in2(_gnd_net_),
            .in3(N__49613),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(elapsed_time_ns_1_RNI57CN9_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_18_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_18_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_18_20_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_18_20_7  (
            .in0(N__49614),
            .in1(_gnd_net_),
            .in2(N__48203),
            .in3(N__48074),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49058),
            .ce(N__50047),
            .sr(N__48580));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_21_0 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_21_0  (
            .in0(N__50144),
            .in1(N__48004),
            .in2(N__50213),
            .in3(N__47989),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_18_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_18_21_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_18_21_1  (
            .in0(N__48168),
            .in1(N__48147),
            .in2(N__48113),
            .in3(N__48066),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_18_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_18_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_18_21_2  (
            .in0(N__48044),
            .in1(N__48035),
            .in2(N__48026),
            .in3(N__47774),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_4 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_4  (
            .in0(N__50143),
            .in1(N__48003),
            .in2(N__50212),
            .in3(N__47988),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_18_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_18_21_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_18_21_6  (
            .in0(N__47913),
            .in1(N__47958),
            .in2(_gnd_net_),
            .in3(N__49593),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_21_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_21_7  (
            .in0(N__47885),
            .in1(N__47844),
            .in2(N__49777),
            .in3(N__47801),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_18_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_18_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_18_22_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_27_LC_18_22_2  (
            .in0(N__50267),
            .in1(N__50237),
            .in2(_gnd_net_),
            .in3(N__49458),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49044),
            .ce(N__49983),
            .sr(N__48596));
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_18_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_18_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_18_22_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_26_LC_18_22_4  (
            .in0(N__50198),
            .in1(N__50173),
            .in2(_gnd_net_),
            .in3(N__49457),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49044),
            .ce(N__49983),
            .sr(N__48596));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_17_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_17_0  (
            .in0(_gnd_net_),
            .in1(N__50135),
            .in2(_gnd_net_),
            .in3(N__50100),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_20_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_20_18_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_20_18_5  (
            .in0(N__49659),
            .in1(N__49713),
            .in2(_gnd_net_),
            .in3(N__49617),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_21_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_21_3  (
            .in0(N__49734),
            .in1(N__49773),
            .in2(_gnd_net_),
            .in3(N__49639),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_20_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_20_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_20_24_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_20_24_2  (
            .in0(N__49715),
            .in1(N__49667),
            .in2(_gnd_net_),
            .in3(N__49555),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49045),
            .ce(N__48721),
            .sr(N__48615));
endmodule // MAIN
