-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 4 2025 00:09:05

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    T01 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__48428\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48380\ : std_logic;
signal \N__48379\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48025\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46718\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46612\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45767\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45703\ : std_logic;
signal \N__45700\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45320\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43788\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42665\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42332\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41906\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41048\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\ : std_logic;
signal \N_38_i_i\ : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_154\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_149\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_153\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_155\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_2_18_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_53\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_3_12_0_\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_62\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_19\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_RNOZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_103_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTIZ0Z1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_434_i\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_30\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \elapsed_time_ns_1_RNI62CED1_0_19_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_315_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_315\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_283_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_307\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIIU2KD1_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIDP2KD1_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_327\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_19\ : std_logic;
signal s3_phy_c : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_72\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\ : std_logic;
signal \elapsed_time_ns_1_RNIL13KD1_0_9_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI1BND11_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI1BND11_0_29_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIT6ND11_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNI0AND11_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNIV8ND11_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNIT6ND11_0_25_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIU7ND11_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNIP2ND11_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNIS5ND11_0_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_17\ : std_logic;
signal \elapsed_time_ns_1_RNIQ3ND11_0_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIR4ND11_0_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\ : std_logic;
signal \elapsed_time_ns_1_RNI3VBED1_0_16_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIA3DJ11_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNI40CED1_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNIA3DJ11_0_4_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI51CED1_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI62CED1_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_328\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_337\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNIQURR91_0_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNINVLD11_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIQ2MD11_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNINVLD11_0_10_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIP1MD11_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_319_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI1TBED1_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_275\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_319\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0Z0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNIQ4OD11_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_278\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \elapsed_time_ns_1_RNID6DJ11_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIE7DJ11_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIB4DJ11_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIS4MD11_0_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_1_sqmuxa\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_1_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_latched2_0\ : std_logic;
signal s4_phy_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_103\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_8\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_382_i_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIP3OD11_0_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_432_i\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNIO0MD11_0_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\ : std_logic;
signal \T01_c\ : std_logic;
signal \T12_c\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_inst2.time_passed_RNI9M3O_cascade_\ : std_logic;
signal \phase_controller_inst2.time_passed_RNI9M3O\ : std_logic;
signal \T23_c\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \T45_c\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_433_i\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \bfn_13_5_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_435_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_1_sqmuxa_cascade_\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_0_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \elapsed_time_ns_1_RNI3VBED1_0_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16\ : std_logic;
signal start_stop_c : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal s2_phy_c : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_359_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_345\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_345_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_341\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_434_i_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_348\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_367\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_349_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_363_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_380\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_378\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_359_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_347\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_347_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_365\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIUDIF91_0_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \phase_controller_inst1.N_55_cascade_\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_latched2_0\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_1_sqmuxa\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_381\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_358\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNI1HIF91_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI0GIF91_0_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \elapsed_time_ns_1_RNI2IIF91_0_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\ : std_logic;
signal \elapsed_time_ns_1_RNIL13KD1_0_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQZ0Z1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_start_latched2_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.N_1609_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal \elapsed_time_ns_1_RNI81DJ11_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_432_i_g\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_382_i\ : std_logic;
signal \elapsed_time_ns_1_RNIO1ND11_0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.timer_s1.N_166_i\ : std_logic;
signal s1_phy_c : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal state_3 : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \elapsed_time_ns_1_RNICG2591_0_4_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_241_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_13\ : std_logic;
signal \elapsed_time_ns_1_RNISAHF91_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNIQ8HF91_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIP7HF91_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIR9HF91_0_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \elapsed_time_ns_1_RNIRAIF91_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNIRBJF91_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNI3JIF91_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNIRAIF91_0_21_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIQ9IF91_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNISBIF91_0_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\ : std_logic;
signal \elapsed_time_ns_1_RNIHI4DM1_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_18\ : std_logic;
signal \elapsed_time_ns_1_RNIGH4DM1_0_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_241\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_9\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.N_56\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_167_i\ : std_logic;
signal \elapsed_time_ns_1_RNIIJ4DM1_0_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_219\ : std_logic;
signal \elapsed_time_ns_1_RNIAE2591_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6\ : std_logic;
signal \elapsed_time_ns_1_RNIGK2591_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_247\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_247_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_251\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\ : std_logic;
signal \elapsed_time_ns_1_RNI1OL2M1_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNIDE4DM1_0_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_244\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNIUCHF91_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_211_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \elapsed_time_ns_1_RNIFG4DM1_0_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1\ : std_logic;
signal \elapsed_time_ns_1_RNIPFL2M1_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_235\ : std_logic;
signal \elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_1\ : std_logic;
signal \elapsed_time_ns_1_RNIUKL2M1_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_5\ : std_logic;
signal \elapsed_time_ns_1_RNIFJ2591_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_7\ : std_logic;
signal \elapsed_time_ns_1_RNICG2591_0_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_4\ : std_logic;
signal \elapsed_time_ns_1_RNISCJF91_0_31\ : std_logic;
signal \elapsed_time_ns_1_RNIDH2591_0_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\ : std_logic;
signal \elapsed_time_ns_1_RNIRHL2M1_0_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_1_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_start_latched2_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8IZ0Z2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input_0_31\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_18_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \current_shift_inst.timer_s1.N_166_i_g\ : std_logic;
signal red_c_g : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal reset_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21356\&\N__21349\&\N__21354\&\N__21348\&\N__21355\&\N__21347\&\N__21357\&\N__21344\&\N__21350\&\N__21343\&\N__21351\&\N__21345\&\N__21352\&\N__21346\&\N__21353\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__39009\&\N__39059\&'0'&'0'&'0'&\N__39057\&\N__39008\&\N__39058\&\N__39007\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21395\&\N__21440\&\N__21396\&\N__21441\&\N__21397\&\N__19998\&\N__20025\&\N__19917\&\N__19956\&\N__20286\&\N__18845\&\N__18825\&\N__18764\&\N__18782\&\N__18797\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__38996\&\N__38993\&'0'&'0'&'0'&\N__38991\&\N__38995\&\N__38992\&\N__38994\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__20615\,
            RESETB => \N__18575\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__39010\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__39056\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__38997\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__38990\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__48426\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48428\,
            DIN => \N__48427\,
            DOUT => \N__48426\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48428\,
            PADOUT => \N__48427\,
            PADIN => \N__48426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48417\,
            DIN => \N__48416\,
            DOUT => \N__48415\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48417\,
            PADOUT => \N__48416\,
            PADIN => \N__48415\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31658\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48408\,
            DIN => \N__48407\,
            DOUT => \N__48406\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48408\,
            PADOUT => \N__48407\,
            PADIN => \N__48406\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48399\,
            DIN => \N__48398\,
            DOUT => \N__48397\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48399\,
            PADOUT => \N__48398\,
            PADIN => \N__48397\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48390\,
            DIN => \N__48389\,
            DOUT => \N__48388\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48390\,
            PADOUT => \N__48389\,
            PADIN => \N__48388\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32039\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48381\,
            DIN => \N__48380\,
            DOUT => \N__48379\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48381\,
            PADOUT => \N__48380\,
            PADIN => \N__48379\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20333\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48372\,
            DIN => \N__48371\,
            DOUT => \N__48370\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48372\,
            PADOUT => \N__48371\,
            PADIN => \N__48370\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48363\,
            DIN => \N__48362\,
            DOUT => \N__48361\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48363\,
            PADOUT => \N__48362\,
            PADIN => \N__48361\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34076\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48354\,
            DIN => \N__48353\,
            DOUT => \N__48352\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48354\,
            PADOUT => \N__48353\,
            PADIN => \N__48352\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32183\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48345\,
            DIN => \N__48344\,
            DOUT => \N__48343\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48345\,
            PADOUT => \N__48344\,
            PADIN => \N__48343\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48336\,
            DIN => \N__48335\,
            DOUT => \N__48334\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48336\,
            PADOUT => \N__48335\,
            PADIN => \N__48334\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__37613\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48327\,
            DIN => \N__48326\,
            DOUT => \N__48325\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48327\,
            PADOUT => \N__48326\,
            PADIN => \N__48325\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27644\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48318\,
            DIN => \N__48317\,
            DOUT => \N__48316\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48318\,
            PADOUT => \N__48317\,
            PADIN => \N__48316\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48309\,
            DIN => \N__48308\,
            DOUT => \N__48307\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48309\,
            PADOUT => \N__48308\,
            PADIN => \N__48307\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25190\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48300\,
            DIN => \N__48299\,
            DOUT => \N__48298\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48300\,
            PADOUT => \N__48299\,
            PADIN => \N__48298\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32348\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48291\,
            DIN => \N__48290\,
            DOUT => \N__48289\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48291\,
            PADOUT => \N__48290\,
            PADIN => \N__48289\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48282\,
            DIN => \N__48281\,
            DOUT => \N__48280\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48282\,
            PADOUT => \N__48281\,
            PADIN => \N__48280\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11474\ : InMux
    port map (
            O => \N__48263\,
            I => \N__48257\
        );

    \I__11473\ : InMux
    port map (
            O => \N__48262\,
            I => \N__48257\
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__48257\,
            I => \N__48253\
        );

    \I__11471\ : InMux
    port map (
            O => \N__48256\,
            I => \N__48250\
        );

    \I__11470\ : Span4Mux_h
    port map (
            O => \N__48253\,
            I => \N__48247\
        );

    \I__11469\ : LocalMux
    port map (
            O => \N__48250\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__11468\ : Odrv4
    port map (
            O => \N__48247\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__11467\ : InMux
    port map (
            O => \N__48242\,
            I => \N__48239\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__48239\,
            I => \N__48234\
        );

    \I__11465\ : InMux
    port map (
            O => \N__48238\,
            I => \N__48231\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48237\,
            I => \N__48228\
        );

    \I__11463\ : Span4Mux_v
    port map (
            O => \N__48234\,
            I => \N__48225\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__48231\,
            I => \N__48220\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__48228\,
            I => \N__48220\
        );

    \I__11460\ : Span4Mux_h
    port map (
            O => \N__48225\,
            I => \N__48214\
        );

    \I__11459\ : Span4Mux_v
    port map (
            O => \N__48220\,
            I => \N__48214\
        );

    \I__11458\ : InMux
    port map (
            O => \N__48219\,
            I => \N__48211\
        );

    \I__11457\ : Odrv4
    port map (
            O => \N__48214\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__48211\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__11455\ : InMux
    port map (
            O => \N__48206\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__11454\ : CascadeMux
    port map (
            O => \N__48203\,
            I => \N__48199\
        );

    \I__11453\ : CascadeMux
    port map (
            O => \N__48202\,
            I => \N__48196\
        );

    \I__11452\ : InMux
    port map (
            O => \N__48199\,
            I => \N__48193\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48196\,
            I => \N__48190\
        );

    \I__11450\ : LocalMux
    port map (
            O => \N__48193\,
            I => \N__48186\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__48190\,
            I => \N__48183\
        );

    \I__11448\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48180\
        );

    \I__11447\ : Span4Mux_h
    port map (
            O => \N__48186\,
            I => \N__48177\
        );

    \I__11446\ : Span4Mux_h
    port map (
            O => \N__48183\,
            I => \N__48174\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__48180\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__11444\ : Odrv4
    port map (
            O => \N__48177\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__11443\ : Odrv4
    port map (
            O => \N__48174\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__11442\ : InMux
    port map (
            O => \N__48167\,
            I => \N__48163\
        );

    \I__11441\ : CascadeMux
    port map (
            O => \N__48166\,
            I => \N__48160\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__48163\,
            I => \N__48156\
        );

    \I__11439\ : InMux
    port map (
            O => \N__48160\,
            I => \N__48153\
        );

    \I__11438\ : CascadeMux
    port map (
            O => \N__48159\,
            I => \N__48150\
        );

    \I__11437\ : Span4Mux_v
    port map (
            O => \N__48156\,
            I => \N__48147\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__48153\,
            I => \N__48144\
        );

    \I__11435\ : InMux
    port map (
            O => \N__48150\,
            I => \N__48141\
        );

    \I__11434\ : Span4Mux_h
    port map (
            O => \N__48147\,
            I => \N__48133\
        );

    \I__11433\ : Span4Mux_v
    port map (
            O => \N__48144\,
            I => \N__48133\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__48141\,
            I => \N__48133\
        );

    \I__11431\ : InMux
    port map (
            O => \N__48140\,
            I => \N__48130\
        );

    \I__11430\ : Odrv4
    port map (
            O => \N__48133\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__48130\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11428\ : InMux
    port map (
            O => \N__48125\,
            I => \bfn_18_22_0_\
        );

    \I__11427\ : CascadeMux
    port map (
            O => \N__48122\,
            I => \N__48118\
        );

    \I__11426\ : CascadeMux
    port map (
            O => \N__48121\,
            I => \N__48115\
        );

    \I__11425\ : InMux
    port map (
            O => \N__48118\,
            I => \N__48112\
        );

    \I__11424\ : InMux
    port map (
            O => \N__48115\,
            I => \N__48109\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__48112\,
            I => \N__48105\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__48109\,
            I => \N__48102\
        );

    \I__11421\ : InMux
    port map (
            O => \N__48108\,
            I => \N__48099\
        );

    \I__11420\ : Span4Mux_h
    port map (
            O => \N__48105\,
            I => \N__48096\
        );

    \I__11419\ : Span4Mux_h
    port map (
            O => \N__48102\,
            I => \N__48093\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__48099\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__11417\ : Odrv4
    port map (
            O => \N__48096\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__11416\ : Odrv4
    port map (
            O => \N__48093\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__11415\ : InMux
    port map (
            O => \N__48086\,
            I => \N__48079\
        );

    \I__11414\ : InMux
    port map (
            O => \N__48085\,
            I => \N__48079\
        );

    \I__11413\ : InMux
    port map (
            O => \N__48084\,
            I => \N__48076\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__48079\,
            I => \N__48073\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__48076\,
            I => \N__48070\
        );

    \I__11410\ : Span4Mux_v
    port map (
            O => \N__48073\,
            I => \N__48067\
        );

    \I__11409\ : Span12Mux_v
    port map (
            O => \N__48070\,
            I => \N__48063\
        );

    \I__11408\ : Span4Mux_v
    port map (
            O => \N__48067\,
            I => \N__48060\
        );

    \I__11407\ : InMux
    port map (
            O => \N__48066\,
            I => \N__48057\
        );

    \I__11406\ : Odrv12
    port map (
            O => \N__48063\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11405\ : Odrv4
    port map (
            O => \N__48060\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48057\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__11403\ : InMux
    port map (
            O => \N__48050\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__11402\ : InMux
    port map (
            O => \N__48047\,
            I => \N__48044\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__48044\,
            I => \N__48040\
        );

    \I__11400\ : InMux
    port map (
            O => \N__48043\,
            I => \N__48037\
        );

    \I__11399\ : Span4Mux_h
    port map (
            O => \N__48040\,
            I => \N__48034\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__48037\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__11397\ : Odrv4
    port map (
            O => \N__48034\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__11396\ : CascadeMux
    port map (
            O => \N__48029\,
            I => \N__48026\
        );

    \I__11395\ : InMux
    port map (
            O => \N__48026\,
            I => \N__48021\
        );

    \I__11394\ : InMux
    port map (
            O => \N__48025\,
            I => \N__48018\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48024\,
            I => \N__48015\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__48021\,
            I => \N__48010\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__48018\,
            I => \N__48010\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__48015\,
            I => \N__48005\
        );

    \I__11389\ : Span4Mux_v
    port map (
            O => \N__48010\,
            I => \N__48005\
        );

    \I__11388\ : Odrv4
    port map (
            O => \N__48005\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__11387\ : InMux
    port map (
            O => \N__48002\,
            I => \N__47998\
        );

    \I__11386\ : InMux
    port map (
            O => \N__48001\,
            I => \N__47995\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__47998\,
            I => \N__47992\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__47995\,
            I => \N__47988\
        );

    \I__11383\ : Span4Mux_v
    port map (
            O => \N__47992\,
            I => \N__47985\
        );

    \I__11382\ : InMux
    port map (
            O => \N__47991\,
            I => \N__47982\
        );

    \I__11381\ : Span12Mux_h
    port map (
            O => \N__47988\,
            I => \N__47978\
        );

    \I__11380\ : Span4Mux_h
    port map (
            O => \N__47985\,
            I => \N__47973\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__47982\,
            I => \N__47973\
        );

    \I__11378\ : InMux
    port map (
            O => \N__47981\,
            I => \N__47970\
        );

    \I__11377\ : Odrv12
    port map (
            O => \N__47978\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__11376\ : Odrv4
    port map (
            O => \N__47973\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__47970\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__11374\ : InMux
    port map (
            O => \N__47963\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__11373\ : InMux
    port map (
            O => \N__47960\,
            I => \N__47957\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__47957\,
            I => \N__47953\
        );

    \I__11371\ : InMux
    port map (
            O => \N__47956\,
            I => \N__47950\
        );

    \I__11370\ : Span4Mux_h
    port map (
            O => \N__47953\,
            I => \N__47947\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__47950\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__11368\ : Odrv4
    port map (
            O => \N__47947\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__11367\ : CascadeMux
    port map (
            O => \N__47942\,
            I => \N__47939\
        );

    \I__11366\ : InMux
    port map (
            O => \N__47939\,
            I => \N__47935\
        );

    \I__11365\ : InMux
    port map (
            O => \N__47938\,
            I => \N__47932\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__47935\,
            I => \N__47926\
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__47932\,
            I => \N__47926\
        );

    \I__11362\ : InMux
    port map (
            O => \N__47931\,
            I => \N__47923\
        );

    \I__11361\ : Span4Mux_v
    port map (
            O => \N__47926\,
            I => \N__47920\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__47923\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__11359\ : Odrv4
    port map (
            O => \N__47920\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__11358\ : InMux
    port map (
            O => \N__47915\,
            I => \N__47911\
        );

    \I__11357\ : InMux
    port map (
            O => \N__47914\,
            I => \N__47908\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__47911\,
            I => \N__47904\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__47908\,
            I => \N__47901\
        );

    \I__11354\ : InMux
    port map (
            O => \N__47907\,
            I => \N__47898\
        );

    \I__11353\ : Span4Mux_v
    port map (
            O => \N__47904\,
            I => \N__47894\
        );

    \I__11352\ : Span4Mux_v
    port map (
            O => \N__47901\,
            I => \N__47889\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__47898\,
            I => \N__47889\
        );

    \I__11350\ : InMux
    port map (
            O => \N__47897\,
            I => \N__47886\
        );

    \I__11349\ : Odrv4
    port map (
            O => \N__47894\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__11348\ : Odrv4
    port map (
            O => \N__47889\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__47886\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__11346\ : InMux
    port map (
            O => \N__47879\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__11345\ : ClkMux
    port map (
            O => \N__47876\,
            I => \N__47519\
        );

    \I__11344\ : ClkMux
    port map (
            O => \N__47875\,
            I => \N__47519\
        );

    \I__11343\ : ClkMux
    port map (
            O => \N__47874\,
            I => \N__47519\
        );

    \I__11342\ : ClkMux
    port map (
            O => \N__47873\,
            I => \N__47519\
        );

    \I__11341\ : ClkMux
    port map (
            O => \N__47872\,
            I => \N__47519\
        );

    \I__11340\ : ClkMux
    port map (
            O => \N__47871\,
            I => \N__47519\
        );

    \I__11339\ : ClkMux
    port map (
            O => \N__47870\,
            I => \N__47519\
        );

    \I__11338\ : ClkMux
    port map (
            O => \N__47869\,
            I => \N__47519\
        );

    \I__11337\ : ClkMux
    port map (
            O => \N__47868\,
            I => \N__47519\
        );

    \I__11336\ : ClkMux
    port map (
            O => \N__47867\,
            I => \N__47519\
        );

    \I__11335\ : ClkMux
    port map (
            O => \N__47866\,
            I => \N__47519\
        );

    \I__11334\ : ClkMux
    port map (
            O => \N__47865\,
            I => \N__47519\
        );

    \I__11333\ : ClkMux
    port map (
            O => \N__47864\,
            I => \N__47519\
        );

    \I__11332\ : ClkMux
    port map (
            O => \N__47863\,
            I => \N__47519\
        );

    \I__11331\ : ClkMux
    port map (
            O => \N__47862\,
            I => \N__47519\
        );

    \I__11330\ : ClkMux
    port map (
            O => \N__47861\,
            I => \N__47519\
        );

    \I__11329\ : ClkMux
    port map (
            O => \N__47860\,
            I => \N__47519\
        );

    \I__11328\ : ClkMux
    port map (
            O => \N__47859\,
            I => \N__47519\
        );

    \I__11327\ : ClkMux
    port map (
            O => \N__47858\,
            I => \N__47519\
        );

    \I__11326\ : ClkMux
    port map (
            O => \N__47857\,
            I => \N__47519\
        );

    \I__11325\ : ClkMux
    port map (
            O => \N__47856\,
            I => \N__47519\
        );

    \I__11324\ : ClkMux
    port map (
            O => \N__47855\,
            I => \N__47519\
        );

    \I__11323\ : ClkMux
    port map (
            O => \N__47854\,
            I => \N__47519\
        );

    \I__11322\ : ClkMux
    port map (
            O => \N__47853\,
            I => \N__47519\
        );

    \I__11321\ : ClkMux
    port map (
            O => \N__47852\,
            I => \N__47519\
        );

    \I__11320\ : ClkMux
    port map (
            O => \N__47851\,
            I => \N__47519\
        );

    \I__11319\ : ClkMux
    port map (
            O => \N__47850\,
            I => \N__47519\
        );

    \I__11318\ : ClkMux
    port map (
            O => \N__47849\,
            I => \N__47519\
        );

    \I__11317\ : ClkMux
    port map (
            O => \N__47848\,
            I => \N__47519\
        );

    \I__11316\ : ClkMux
    port map (
            O => \N__47847\,
            I => \N__47519\
        );

    \I__11315\ : ClkMux
    port map (
            O => \N__47846\,
            I => \N__47519\
        );

    \I__11314\ : ClkMux
    port map (
            O => \N__47845\,
            I => \N__47519\
        );

    \I__11313\ : ClkMux
    port map (
            O => \N__47844\,
            I => \N__47519\
        );

    \I__11312\ : ClkMux
    port map (
            O => \N__47843\,
            I => \N__47519\
        );

    \I__11311\ : ClkMux
    port map (
            O => \N__47842\,
            I => \N__47519\
        );

    \I__11310\ : ClkMux
    port map (
            O => \N__47841\,
            I => \N__47519\
        );

    \I__11309\ : ClkMux
    port map (
            O => \N__47840\,
            I => \N__47519\
        );

    \I__11308\ : ClkMux
    port map (
            O => \N__47839\,
            I => \N__47519\
        );

    \I__11307\ : ClkMux
    port map (
            O => \N__47838\,
            I => \N__47519\
        );

    \I__11306\ : ClkMux
    port map (
            O => \N__47837\,
            I => \N__47519\
        );

    \I__11305\ : ClkMux
    port map (
            O => \N__47836\,
            I => \N__47519\
        );

    \I__11304\ : ClkMux
    port map (
            O => \N__47835\,
            I => \N__47519\
        );

    \I__11303\ : ClkMux
    port map (
            O => \N__47834\,
            I => \N__47519\
        );

    \I__11302\ : ClkMux
    port map (
            O => \N__47833\,
            I => \N__47519\
        );

    \I__11301\ : ClkMux
    port map (
            O => \N__47832\,
            I => \N__47519\
        );

    \I__11300\ : ClkMux
    port map (
            O => \N__47831\,
            I => \N__47519\
        );

    \I__11299\ : ClkMux
    port map (
            O => \N__47830\,
            I => \N__47519\
        );

    \I__11298\ : ClkMux
    port map (
            O => \N__47829\,
            I => \N__47519\
        );

    \I__11297\ : ClkMux
    port map (
            O => \N__47828\,
            I => \N__47519\
        );

    \I__11296\ : ClkMux
    port map (
            O => \N__47827\,
            I => \N__47519\
        );

    \I__11295\ : ClkMux
    port map (
            O => \N__47826\,
            I => \N__47519\
        );

    \I__11294\ : ClkMux
    port map (
            O => \N__47825\,
            I => \N__47519\
        );

    \I__11293\ : ClkMux
    port map (
            O => \N__47824\,
            I => \N__47519\
        );

    \I__11292\ : ClkMux
    port map (
            O => \N__47823\,
            I => \N__47519\
        );

    \I__11291\ : ClkMux
    port map (
            O => \N__47822\,
            I => \N__47519\
        );

    \I__11290\ : ClkMux
    port map (
            O => \N__47821\,
            I => \N__47519\
        );

    \I__11289\ : ClkMux
    port map (
            O => \N__47820\,
            I => \N__47519\
        );

    \I__11288\ : ClkMux
    port map (
            O => \N__47819\,
            I => \N__47519\
        );

    \I__11287\ : ClkMux
    port map (
            O => \N__47818\,
            I => \N__47519\
        );

    \I__11286\ : ClkMux
    port map (
            O => \N__47817\,
            I => \N__47519\
        );

    \I__11285\ : ClkMux
    port map (
            O => \N__47816\,
            I => \N__47519\
        );

    \I__11284\ : ClkMux
    port map (
            O => \N__47815\,
            I => \N__47519\
        );

    \I__11283\ : ClkMux
    port map (
            O => \N__47814\,
            I => \N__47519\
        );

    \I__11282\ : ClkMux
    port map (
            O => \N__47813\,
            I => \N__47519\
        );

    \I__11281\ : ClkMux
    port map (
            O => \N__47812\,
            I => \N__47519\
        );

    \I__11280\ : ClkMux
    port map (
            O => \N__47811\,
            I => \N__47519\
        );

    \I__11279\ : ClkMux
    port map (
            O => \N__47810\,
            I => \N__47519\
        );

    \I__11278\ : ClkMux
    port map (
            O => \N__47809\,
            I => \N__47519\
        );

    \I__11277\ : ClkMux
    port map (
            O => \N__47808\,
            I => \N__47519\
        );

    \I__11276\ : ClkMux
    port map (
            O => \N__47807\,
            I => \N__47519\
        );

    \I__11275\ : ClkMux
    port map (
            O => \N__47806\,
            I => \N__47519\
        );

    \I__11274\ : ClkMux
    port map (
            O => \N__47805\,
            I => \N__47519\
        );

    \I__11273\ : ClkMux
    port map (
            O => \N__47804\,
            I => \N__47519\
        );

    \I__11272\ : ClkMux
    port map (
            O => \N__47803\,
            I => \N__47519\
        );

    \I__11271\ : ClkMux
    port map (
            O => \N__47802\,
            I => \N__47519\
        );

    \I__11270\ : ClkMux
    port map (
            O => \N__47801\,
            I => \N__47519\
        );

    \I__11269\ : ClkMux
    port map (
            O => \N__47800\,
            I => \N__47519\
        );

    \I__11268\ : ClkMux
    port map (
            O => \N__47799\,
            I => \N__47519\
        );

    \I__11267\ : ClkMux
    port map (
            O => \N__47798\,
            I => \N__47519\
        );

    \I__11266\ : ClkMux
    port map (
            O => \N__47797\,
            I => \N__47519\
        );

    \I__11265\ : ClkMux
    port map (
            O => \N__47796\,
            I => \N__47519\
        );

    \I__11264\ : ClkMux
    port map (
            O => \N__47795\,
            I => \N__47519\
        );

    \I__11263\ : ClkMux
    port map (
            O => \N__47794\,
            I => \N__47519\
        );

    \I__11262\ : ClkMux
    port map (
            O => \N__47793\,
            I => \N__47519\
        );

    \I__11261\ : ClkMux
    port map (
            O => \N__47792\,
            I => \N__47519\
        );

    \I__11260\ : ClkMux
    port map (
            O => \N__47791\,
            I => \N__47519\
        );

    \I__11259\ : ClkMux
    port map (
            O => \N__47790\,
            I => \N__47519\
        );

    \I__11258\ : ClkMux
    port map (
            O => \N__47789\,
            I => \N__47519\
        );

    \I__11257\ : ClkMux
    port map (
            O => \N__47788\,
            I => \N__47519\
        );

    \I__11256\ : ClkMux
    port map (
            O => \N__47787\,
            I => \N__47519\
        );

    \I__11255\ : ClkMux
    port map (
            O => \N__47786\,
            I => \N__47519\
        );

    \I__11254\ : ClkMux
    port map (
            O => \N__47785\,
            I => \N__47519\
        );

    \I__11253\ : ClkMux
    port map (
            O => \N__47784\,
            I => \N__47519\
        );

    \I__11252\ : ClkMux
    port map (
            O => \N__47783\,
            I => \N__47519\
        );

    \I__11251\ : ClkMux
    port map (
            O => \N__47782\,
            I => \N__47519\
        );

    \I__11250\ : ClkMux
    port map (
            O => \N__47781\,
            I => \N__47519\
        );

    \I__11249\ : ClkMux
    port map (
            O => \N__47780\,
            I => \N__47519\
        );

    \I__11248\ : ClkMux
    port map (
            O => \N__47779\,
            I => \N__47519\
        );

    \I__11247\ : ClkMux
    port map (
            O => \N__47778\,
            I => \N__47519\
        );

    \I__11246\ : ClkMux
    port map (
            O => \N__47777\,
            I => \N__47519\
        );

    \I__11245\ : ClkMux
    port map (
            O => \N__47776\,
            I => \N__47519\
        );

    \I__11244\ : ClkMux
    port map (
            O => \N__47775\,
            I => \N__47519\
        );

    \I__11243\ : ClkMux
    port map (
            O => \N__47774\,
            I => \N__47519\
        );

    \I__11242\ : ClkMux
    port map (
            O => \N__47773\,
            I => \N__47519\
        );

    \I__11241\ : ClkMux
    port map (
            O => \N__47772\,
            I => \N__47519\
        );

    \I__11240\ : ClkMux
    port map (
            O => \N__47771\,
            I => \N__47519\
        );

    \I__11239\ : ClkMux
    port map (
            O => \N__47770\,
            I => \N__47519\
        );

    \I__11238\ : ClkMux
    port map (
            O => \N__47769\,
            I => \N__47519\
        );

    \I__11237\ : ClkMux
    port map (
            O => \N__47768\,
            I => \N__47519\
        );

    \I__11236\ : ClkMux
    port map (
            O => \N__47767\,
            I => \N__47519\
        );

    \I__11235\ : ClkMux
    port map (
            O => \N__47766\,
            I => \N__47519\
        );

    \I__11234\ : ClkMux
    port map (
            O => \N__47765\,
            I => \N__47519\
        );

    \I__11233\ : ClkMux
    port map (
            O => \N__47764\,
            I => \N__47519\
        );

    \I__11232\ : ClkMux
    port map (
            O => \N__47763\,
            I => \N__47519\
        );

    \I__11231\ : ClkMux
    port map (
            O => \N__47762\,
            I => \N__47519\
        );

    \I__11230\ : ClkMux
    port map (
            O => \N__47761\,
            I => \N__47519\
        );

    \I__11229\ : ClkMux
    port map (
            O => \N__47760\,
            I => \N__47519\
        );

    \I__11228\ : ClkMux
    port map (
            O => \N__47759\,
            I => \N__47519\
        );

    \I__11227\ : ClkMux
    port map (
            O => \N__47758\,
            I => \N__47519\
        );

    \I__11226\ : GlobalMux
    port map (
            O => \N__47519\,
            I => clk_100mhz_0
        );

    \I__11225\ : CEMux
    port map (
            O => \N__47516\,
            I => \N__47489\
        );

    \I__11224\ : CEMux
    port map (
            O => \N__47515\,
            I => \N__47489\
        );

    \I__11223\ : CEMux
    port map (
            O => \N__47514\,
            I => \N__47489\
        );

    \I__11222\ : CEMux
    port map (
            O => \N__47513\,
            I => \N__47489\
        );

    \I__11221\ : CEMux
    port map (
            O => \N__47512\,
            I => \N__47489\
        );

    \I__11220\ : CEMux
    port map (
            O => \N__47511\,
            I => \N__47489\
        );

    \I__11219\ : CEMux
    port map (
            O => \N__47510\,
            I => \N__47489\
        );

    \I__11218\ : CEMux
    port map (
            O => \N__47509\,
            I => \N__47489\
        );

    \I__11217\ : CEMux
    port map (
            O => \N__47508\,
            I => \N__47489\
        );

    \I__11216\ : GlobalMux
    port map (
            O => \N__47489\,
            I => \N__47486\
        );

    \I__11215\ : gio2CtrlBuf
    port map (
            O => \N__47486\,
            I => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \I__11214\ : InMux
    port map (
            O => \N__47483\,
            I => \N__47466\
        );

    \I__11213\ : InMux
    port map (
            O => \N__47482\,
            I => \N__47463\
        );

    \I__11212\ : InMux
    port map (
            O => \N__47481\,
            I => \N__47460\
        );

    \I__11211\ : InMux
    port map (
            O => \N__47480\,
            I => \N__47457\
        );

    \I__11210\ : InMux
    port map (
            O => \N__47479\,
            I => \N__47454\
        );

    \I__11209\ : InMux
    port map (
            O => \N__47478\,
            I => \N__47449\
        );

    \I__11208\ : InMux
    port map (
            O => \N__47477\,
            I => \N__47449\
        );

    \I__11207\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47444\
        );

    \I__11206\ : InMux
    port map (
            O => \N__47475\,
            I => \N__47444\
        );

    \I__11205\ : InMux
    port map (
            O => \N__47474\,
            I => \N__47439\
        );

    \I__11204\ : InMux
    port map (
            O => \N__47473\,
            I => \N__47439\
        );

    \I__11203\ : InMux
    port map (
            O => \N__47472\,
            I => \N__47434\
        );

    \I__11202\ : InMux
    port map (
            O => \N__47471\,
            I => \N__47434\
        );

    \I__11201\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47431\
        );

    \I__11200\ : InMux
    port map (
            O => \N__47469\,
            I => \N__47428\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__47466\,
            I => \N__47425\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__47463\,
            I => \N__47422\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__47460\,
            I => \N__47419\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__47457\,
            I => \N__47411\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__47454\,
            I => \N__47355\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__47449\,
            I => \N__47346\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__47444\,
            I => \N__47343\
        );

    \I__11192\ : LocalMux
    port map (
            O => \N__47439\,
            I => \N__47336\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__47434\,
            I => \N__47308\
        );

    \I__11190\ : LocalMux
    port map (
            O => \N__47431\,
            I => \N__47296\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__47428\,
            I => \N__47290\
        );

    \I__11188\ : Glb2LocalMux
    port map (
            O => \N__47425\,
            I => \N__47030\
        );

    \I__11187\ : Glb2LocalMux
    port map (
            O => \N__47422\,
            I => \N__47030\
        );

    \I__11186\ : Glb2LocalMux
    port map (
            O => \N__47419\,
            I => \N__47030\
        );

    \I__11185\ : SRMux
    port map (
            O => \N__47418\,
            I => \N__47030\
        );

    \I__11184\ : SRMux
    port map (
            O => \N__47417\,
            I => \N__47030\
        );

    \I__11183\ : SRMux
    port map (
            O => \N__47416\,
            I => \N__47030\
        );

    \I__11182\ : SRMux
    port map (
            O => \N__47415\,
            I => \N__47030\
        );

    \I__11181\ : SRMux
    port map (
            O => \N__47414\,
            I => \N__47030\
        );

    \I__11180\ : Glb2LocalMux
    port map (
            O => \N__47411\,
            I => \N__47030\
        );

    \I__11179\ : SRMux
    port map (
            O => \N__47410\,
            I => \N__47030\
        );

    \I__11178\ : SRMux
    port map (
            O => \N__47409\,
            I => \N__47030\
        );

    \I__11177\ : SRMux
    port map (
            O => \N__47408\,
            I => \N__47030\
        );

    \I__11176\ : SRMux
    port map (
            O => \N__47407\,
            I => \N__47030\
        );

    \I__11175\ : SRMux
    port map (
            O => \N__47406\,
            I => \N__47030\
        );

    \I__11174\ : SRMux
    port map (
            O => \N__47405\,
            I => \N__47030\
        );

    \I__11173\ : SRMux
    port map (
            O => \N__47404\,
            I => \N__47030\
        );

    \I__11172\ : SRMux
    port map (
            O => \N__47403\,
            I => \N__47030\
        );

    \I__11171\ : SRMux
    port map (
            O => \N__47402\,
            I => \N__47030\
        );

    \I__11170\ : SRMux
    port map (
            O => \N__47401\,
            I => \N__47030\
        );

    \I__11169\ : SRMux
    port map (
            O => \N__47400\,
            I => \N__47030\
        );

    \I__11168\ : SRMux
    port map (
            O => \N__47399\,
            I => \N__47030\
        );

    \I__11167\ : SRMux
    port map (
            O => \N__47398\,
            I => \N__47030\
        );

    \I__11166\ : SRMux
    port map (
            O => \N__47397\,
            I => \N__47030\
        );

    \I__11165\ : SRMux
    port map (
            O => \N__47396\,
            I => \N__47030\
        );

    \I__11164\ : SRMux
    port map (
            O => \N__47395\,
            I => \N__47030\
        );

    \I__11163\ : SRMux
    port map (
            O => \N__47394\,
            I => \N__47030\
        );

    \I__11162\ : SRMux
    port map (
            O => \N__47393\,
            I => \N__47030\
        );

    \I__11161\ : SRMux
    port map (
            O => \N__47392\,
            I => \N__47030\
        );

    \I__11160\ : SRMux
    port map (
            O => \N__47391\,
            I => \N__47030\
        );

    \I__11159\ : SRMux
    port map (
            O => \N__47390\,
            I => \N__47030\
        );

    \I__11158\ : SRMux
    port map (
            O => \N__47389\,
            I => \N__47030\
        );

    \I__11157\ : SRMux
    port map (
            O => \N__47388\,
            I => \N__47030\
        );

    \I__11156\ : SRMux
    port map (
            O => \N__47387\,
            I => \N__47030\
        );

    \I__11155\ : SRMux
    port map (
            O => \N__47386\,
            I => \N__47030\
        );

    \I__11154\ : SRMux
    port map (
            O => \N__47385\,
            I => \N__47030\
        );

    \I__11153\ : SRMux
    port map (
            O => \N__47384\,
            I => \N__47030\
        );

    \I__11152\ : SRMux
    port map (
            O => \N__47383\,
            I => \N__47030\
        );

    \I__11151\ : SRMux
    port map (
            O => \N__47382\,
            I => \N__47030\
        );

    \I__11150\ : SRMux
    port map (
            O => \N__47381\,
            I => \N__47030\
        );

    \I__11149\ : SRMux
    port map (
            O => \N__47380\,
            I => \N__47030\
        );

    \I__11148\ : SRMux
    port map (
            O => \N__47379\,
            I => \N__47030\
        );

    \I__11147\ : SRMux
    port map (
            O => \N__47378\,
            I => \N__47030\
        );

    \I__11146\ : SRMux
    port map (
            O => \N__47377\,
            I => \N__47030\
        );

    \I__11145\ : SRMux
    port map (
            O => \N__47376\,
            I => \N__47030\
        );

    \I__11144\ : SRMux
    port map (
            O => \N__47375\,
            I => \N__47030\
        );

    \I__11143\ : SRMux
    port map (
            O => \N__47374\,
            I => \N__47030\
        );

    \I__11142\ : SRMux
    port map (
            O => \N__47373\,
            I => \N__47030\
        );

    \I__11141\ : SRMux
    port map (
            O => \N__47372\,
            I => \N__47030\
        );

    \I__11140\ : SRMux
    port map (
            O => \N__47371\,
            I => \N__47030\
        );

    \I__11139\ : SRMux
    port map (
            O => \N__47370\,
            I => \N__47030\
        );

    \I__11138\ : SRMux
    port map (
            O => \N__47369\,
            I => \N__47030\
        );

    \I__11137\ : SRMux
    port map (
            O => \N__47368\,
            I => \N__47030\
        );

    \I__11136\ : SRMux
    port map (
            O => \N__47367\,
            I => \N__47030\
        );

    \I__11135\ : SRMux
    port map (
            O => \N__47366\,
            I => \N__47030\
        );

    \I__11134\ : SRMux
    port map (
            O => \N__47365\,
            I => \N__47030\
        );

    \I__11133\ : SRMux
    port map (
            O => \N__47364\,
            I => \N__47030\
        );

    \I__11132\ : SRMux
    port map (
            O => \N__47363\,
            I => \N__47030\
        );

    \I__11131\ : SRMux
    port map (
            O => \N__47362\,
            I => \N__47030\
        );

    \I__11130\ : SRMux
    port map (
            O => \N__47361\,
            I => \N__47030\
        );

    \I__11129\ : SRMux
    port map (
            O => \N__47360\,
            I => \N__47030\
        );

    \I__11128\ : SRMux
    port map (
            O => \N__47359\,
            I => \N__47030\
        );

    \I__11127\ : SRMux
    port map (
            O => \N__47358\,
            I => \N__47030\
        );

    \I__11126\ : Glb2LocalMux
    port map (
            O => \N__47355\,
            I => \N__47030\
        );

    \I__11125\ : SRMux
    port map (
            O => \N__47354\,
            I => \N__47030\
        );

    \I__11124\ : SRMux
    port map (
            O => \N__47353\,
            I => \N__47030\
        );

    \I__11123\ : SRMux
    port map (
            O => \N__47352\,
            I => \N__47030\
        );

    \I__11122\ : SRMux
    port map (
            O => \N__47351\,
            I => \N__47030\
        );

    \I__11121\ : SRMux
    port map (
            O => \N__47350\,
            I => \N__47030\
        );

    \I__11120\ : SRMux
    port map (
            O => \N__47349\,
            I => \N__47030\
        );

    \I__11119\ : Glb2LocalMux
    port map (
            O => \N__47346\,
            I => \N__47030\
        );

    \I__11118\ : Glb2LocalMux
    port map (
            O => \N__47343\,
            I => \N__47030\
        );

    \I__11117\ : SRMux
    port map (
            O => \N__47342\,
            I => \N__47030\
        );

    \I__11116\ : SRMux
    port map (
            O => \N__47341\,
            I => \N__47030\
        );

    \I__11115\ : SRMux
    port map (
            O => \N__47340\,
            I => \N__47030\
        );

    \I__11114\ : SRMux
    port map (
            O => \N__47339\,
            I => \N__47030\
        );

    \I__11113\ : Glb2LocalMux
    port map (
            O => \N__47336\,
            I => \N__47030\
        );

    \I__11112\ : SRMux
    port map (
            O => \N__47335\,
            I => \N__47030\
        );

    \I__11111\ : SRMux
    port map (
            O => \N__47334\,
            I => \N__47030\
        );

    \I__11110\ : SRMux
    port map (
            O => \N__47333\,
            I => \N__47030\
        );

    \I__11109\ : SRMux
    port map (
            O => \N__47332\,
            I => \N__47030\
        );

    \I__11108\ : SRMux
    port map (
            O => \N__47331\,
            I => \N__47030\
        );

    \I__11107\ : SRMux
    port map (
            O => \N__47330\,
            I => \N__47030\
        );

    \I__11106\ : SRMux
    port map (
            O => \N__47329\,
            I => \N__47030\
        );

    \I__11105\ : SRMux
    port map (
            O => \N__47328\,
            I => \N__47030\
        );

    \I__11104\ : SRMux
    port map (
            O => \N__47327\,
            I => \N__47030\
        );

    \I__11103\ : SRMux
    port map (
            O => \N__47326\,
            I => \N__47030\
        );

    \I__11102\ : SRMux
    port map (
            O => \N__47325\,
            I => \N__47030\
        );

    \I__11101\ : SRMux
    port map (
            O => \N__47324\,
            I => \N__47030\
        );

    \I__11100\ : SRMux
    port map (
            O => \N__47323\,
            I => \N__47030\
        );

    \I__11099\ : SRMux
    port map (
            O => \N__47322\,
            I => \N__47030\
        );

    \I__11098\ : SRMux
    port map (
            O => \N__47321\,
            I => \N__47030\
        );

    \I__11097\ : SRMux
    port map (
            O => \N__47320\,
            I => \N__47030\
        );

    \I__11096\ : SRMux
    port map (
            O => \N__47319\,
            I => \N__47030\
        );

    \I__11095\ : SRMux
    port map (
            O => \N__47318\,
            I => \N__47030\
        );

    \I__11094\ : SRMux
    port map (
            O => \N__47317\,
            I => \N__47030\
        );

    \I__11093\ : SRMux
    port map (
            O => \N__47316\,
            I => \N__47030\
        );

    \I__11092\ : SRMux
    port map (
            O => \N__47315\,
            I => \N__47030\
        );

    \I__11091\ : SRMux
    port map (
            O => \N__47314\,
            I => \N__47030\
        );

    \I__11090\ : SRMux
    port map (
            O => \N__47313\,
            I => \N__47030\
        );

    \I__11089\ : SRMux
    port map (
            O => \N__47312\,
            I => \N__47030\
        );

    \I__11088\ : SRMux
    port map (
            O => \N__47311\,
            I => \N__47030\
        );

    \I__11087\ : Glb2LocalMux
    port map (
            O => \N__47308\,
            I => \N__47030\
        );

    \I__11086\ : SRMux
    port map (
            O => \N__47307\,
            I => \N__47030\
        );

    \I__11085\ : SRMux
    port map (
            O => \N__47306\,
            I => \N__47030\
        );

    \I__11084\ : SRMux
    port map (
            O => \N__47305\,
            I => \N__47030\
        );

    \I__11083\ : SRMux
    port map (
            O => \N__47304\,
            I => \N__47030\
        );

    \I__11082\ : SRMux
    port map (
            O => \N__47303\,
            I => \N__47030\
        );

    \I__11081\ : SRMux
    port map (
            O => \N__47302\,
            I => \N__47030\
        );

    \I__11080\ : SRMux
    port map (
            O => \N__47301\,
            I => \N__47030\
        );

    \I__11079\ : SRMux
    port map (
            O => \N__47300\,
            I => \N__47030\
        );

    \I__11078\ : SRMux
    port map (
            O => \N__47299\,
            I => \N__47030\
        );

    \I__11077\ : Glb2LocalMux
    port map (
            O => \N__47296\,
            I => \N__47030\
        );

    \I__11076\ : SRMux
    port map (
            O => \N__47295\,
            I => \N__47030\
        );

    \I__11075\ : SRMux
    port map (
            O => \N__47294\,
            I => \N__47030\
        );

    \I__11074\ : SRMux
    port map (
            O => \N__47293\,
            I => \N__47030\
        );

    \I__11073\ : Glb2LocalMux
    port map (
            O => \N__47290\,
            I => \N__47030\
        );

    \I__11072\ : SRMux
    port map (
            O => \N__47289\,
            I => \N__47030\
        );

    \I__11071\ : SRMux
    port map (
            O => \N__47288\,
            I => \N__47030\
        );

    \I__11070\ : SRMux
    port map (
            O => \N__47287\,
            I => \N__47030\
        );

    \I__11069\ : SRMux
    port map (
            O => \N__47286\,
            I => \N__47030\
        );

    \I__11068\ : SRMux
    port map (
            O => \N__47285\,
            I => \N__47030\
        );

    \I__11067\ : SRMux
    port map (
            O => \N__47284\,
            I => \N__47030\
        );

    \I__11066\ : SRMux
    port map (
            O => \N__47283\,
            I => \N__47030\
        );

    \I__11065\ : SRMux
    port map (
            O => \N__47282\,
            I => \N__47030\
        );

    \I__11064\ : SRMux
    port map (
            O => \N__47281\,
            I => \N__47030\
        );

    \I__11063\ : GlobalMux
    port map (
            O => \N__47030\,
            I => \N__47027\
        );

    \I__11062\ : gio2CtrlBuf
    port map (
            O => \N__47027\,
            I => red_c_g
        );

    \I__11061\ : InMux
    port map (
            O => \N__47024\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__11060\ : InMux
    port map (
            O => \N__47021\,
            I => \N__47016\
        );

    \I__11059\ : InMux
    port map (
            O => \N__47020\,
            I => \N__47013\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47019\,
            I => \N__47010\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__47016\,
            I => \N__47007\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__47013\,
            I => \N__47004\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__47010\,
            I => \N__47001\
        );

    \I__11054\ : Span4Mux_v
    port map (
            O => \N__47007\,
            I => \N__46998\
        );

    \I__11053\ : Span4Mux_h
    port map (
            O => \N__47004\,
            I => \N__46995\
        );

    \I__11052\ : Sp12to4
    port map (
            O => \N__47001\,
            I => \N__46992\
        );

    \I__11051\ : Span4Mux_h
    port map (
            O => \N__46998\,
            I => \N__46987\
        );

    \I__11050\ : Span4Mux_h
    port map (
            O => \N__46995\,
            I => \N__46987\
        );

    \I__11049\ : Odrv12
    port map (
            O => \N__46992\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__11048\ : Odrv4
    port map (
            O => \N__46987\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__11047\ : CascadeMux
    port map (
            O => \N__46982\,
            I => \N__46978\
        );

    \I__11046\ : CascadeMux
    port map (
            O => \N__46981\,
            I => \N__46975\
        );

    \I__11045\ : InMux
    port map (
            O => \N__46978\,
            I => \N__46972\
        );

    \I__11044\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46969\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__46972\,
            I => \N__46965\
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__46969\,
            I => \N__46962\
        );

    \I__11041\ : InMux
    port map (
            O => \N__46968\,
            I => \N__46959\
        );

    \I__11040\ : Span4Mux_h
    port map (
            O => \N__46965\,
            I => \N__46956\
        );

    \I__11039\ : Span4Mux_h
    port map (
            O => \N__46962\,
            I => \N__46953\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__46959\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__11037\ : Odrv4
    port map (
            O => \N__46956\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__11036\ : Odrv4
    port map (
            O => \N__46953\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__11035\ : InMux
    port map (
            O => \N__46946\,
            I => \N__46942\
        );

    \I__11034\ : InMux
    port map (
            O => \N__46945\,
            I => \N__46939\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__46942\,
            I => \N__46936\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__46939\,
            I => \N__46930\
        );

    \I__11031\ : Span4Mux_h
    port map (
            O => \N__46936\,
            I => \N__46930\
        );

    \I__11030\ : InMux
    port map (
            O => \N__46935\,
            I => \N__46926\
        );

    \I__11029\ : Span4Mux_h
    port map (
            O => \N__46930\,
            I => \N__46923\
        );

    \I__11028\ : InMux
    port map (
            O => \N__46929\,
            I => \N__46920\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__46926\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__11026\ : Odrv4
    port map (
            O => \N__46923\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__46920\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__11024\ : InMux
    port map (
            O => \N__46913\,
            I => \bfn_18_21_0_\
        );

    \I__11023\ : CascadeMux
    port map (
            O => \N__46910\,
            I => \N__46906\
        );

    \I__11022\ : CascadeMux
    port map (
            O => \N__46909\,
            I => \N__46903\
        );

    \I__11021\ : InMux
    port map (
            O => \N__46906\,
            I => \N__46900\
        );

    \I__11020\ : InMux
    port map (
            O => \N__46903\,
            I => \N__46897\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__46900\,
            I => \N__46893\
        );

    \I__11018\ : LocalMux
    port map (
            O => \N__46897\,
            I => \N__46890\
        );

    \I__11017\ : InMux
    port map (
            O => \N__46896\,
            I => \N__46887\
        );

    \I__11016\ : Span4Mux_h
    port map (
            O => \N__46893\,
            I => \N__46884\
        );

    \I__11015\ : Span4Mux_h
    port map (
            O => \N__46890\,
            I => \N__46881\
        );

    \I__11014\ : LocalMux
    port map (
            O => \N__46887\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__11013\ : Odrv4
    port map (
            O => \N__46884\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__11012\ : Odrv4
    port map (
            O => \N__46881\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__11011\ : InMux
    port map (
            O => \N__46874\,
            I => \N__46869\
        );

    \I__11010\ : InMux
    port map (
            O => \N__46873\,
            I => \N__46864\
        );

    \I__11009\ : InMux
    port map (
            O => \N__46872\,
            I => \N__46864\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__46869\,
            I => \N__46859\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__46864\,
            I => \N__46859\
        );

    \I__11006\ : Span12Mux_v
    port map (
            O => \N__46859\,
            I => \N__46855\
        );

    \I__11005\ : InMux
    port map (
            O => \N__46858\,
            I => \N__46852\
        );

    \I__11004\ : Odrv12
    port map (
            O => \N__46855\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__46852\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__11002\ : InMux
    port map (
            O => \N__46847\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__11001\ : CascadeMux
    port map (
            O => \N__46844\,
            I => \N__46841\
        );

    \I__11000\ : InMux
    port map (
            O => \N__46841\,
            I => \N__46836\
        );

    \I__10999\ : InMux
    port map (
            O => \N__46840\,
            I => \N__46833\
        );

    \I__10998\ : InMux
    port map (
            O => \N__46839\,
            I => \N__46830\
        );

    \I__10997\ : LocalMux
    port map (
            O => \N__46836\,
            I => \N__46825\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__46833\,
            I => \N__46825\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__46830\,
            I => \N__46820\
        );

    \I__10994\ : Span4Mux_v
    port map (
            O => \N__46825\,
            I => \N__46820\
        );

    \I__10993\ : Odrv4
    port map (
            O => \N__46820\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__10992\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46814\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__46814\,
            I => \N__46809\
        );

    \I__10990\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46806\
        );

    \I__10989\ : InMux
    port map (
            O => \N__46812\,
            I => \N__46802\
        );

    \I__10988\ : Span4Mux_v
    port map (
            O => \N__46809\,
            I => \N__46797\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__46806\,
            I => \N__46797\
        );

    \I__10986\ : InMux
    port map (
            O => \N__46805\,
            I => \N__46794\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__46802\,
            I => \N__46791\
        );

    \I__10984\ : Span4Mux_v
    port map (
            O => \N__46797\,
            I => \N__46788\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__46794\,
            I => \N__46785\
        );

    \I__10982\ : Span4Mux_v
    port map (
            O => \N__46791\,
            I => \N__46782\
        );

    \I__10981\ : Odrv4
    port map (
            O => \N__46788\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10980\ : Odrv4
    port map (
            O => \N__46785\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10979\ : Odrv4
    port map (
            O => \N__46782\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10978\ : InMux
    port map (
            O => \N__46775\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__10977\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46766\
        );

    \I__10976\ : InMux
    port map (
            O => \N__46771\,
            I => \N__46766\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__46766\,
            I => \N__46762\
        );

    \I__10974\ : InMux
    port map (
            O => \N__46765\,
            I => \N__46759\
        );

    \I__10973\ : Span4Mux_v
    port map (
            O => \N__46762\,
            I => \N__46756\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__46759\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__10971\ : Odrv4
    port map (
            O => \N__46756\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__10970\ : InMux
    port map (
            O => \N__46751\,
            I => \N__46742\
        );

    \I__10969\ : InMux
    port map (
            O => \N__46750\,
            I => \N__46742\
        );

    \I__10968\ : InMux
    port map (
            O => \N__46749\,
            I => \N__46742\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__46742\,
            I => \N__46739\
        );

    \I__10966\ : Span4Mux_v
    port map (
            O => \N__46739\,
            I => \N__46736\
        );

    \I__10965\ : Span4Mux_h
    port map (
            O => \N__46736\,
            I => \N__46732\
        );

    \I__10964\ : InMux
    port map (
            O => \N__46735\,
            I => \N__46729\
        );

    \I__10963\ : Odrv4
    port map (
            O => \N__46732\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__46729\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__10961\ : InMux
    port map (
            O => \N__46724\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__10960\ : CascadeMux
    port map (
            O => \N__46721\,
            I => \N__46718\
        );

    \I__10959\ : InMux
    port map (
            O => \N__46718\,
            I => \N__46714\
        );

    \I__10958\ : InMux
    port map (
            O => \N__46717\,
            I => \N__46711\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__46714\,
            I => \N__46705\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__46711\,
            I => \N__46705\
        );

    \I__10955\ : InMux
    port map (
            O => \N__46710\,
            I => \N__46702\
        );

    \I__10954\ : Span4Mux_h
    port map (
            O => \N__46705\,
            I => \N__46699\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__46702\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__10952\ : Odrv4
    port map (
            O => \N__46699\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__10951\ : InMux
    port map (
            O => \N__46694\,
            I => \N__46689\
        );

    \I__10950\ : InMux
    port map (
            O => \N__46693\,
            I => \N__46686\
        );

    \I__10949\ : InMux
    port map (
            O => \N__46692\,
            I => \N__46683\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__46689\,
            I => \N__46677\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__46686\,
            I => \N__46677\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__46683\,
            I => \N__46674\
        );

    \I__10945\ : InMux
    port map (
            O => \N__46682\,
            I => \N__46671\
        );

    \I__10944\ : Span4Mux_h
    port map (
            O => \N__46677\,
            I => \N__46668\
        );

    \I__10943\ : Span4Mux_h
    port map (
            O => \N__46674\,
            I => \N__46663\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__46671\,
            I => \N__46663\
        );

    \I__10941\ : Odrv4
    port map (
            O => \N__46668\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10940\ : Odrv4
    port map (
            O => \N__46663\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10939\ : InMux
    port map (
            O => \N__46658\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__10938\ : CascadeMux
    port map (
            O => \N__46655\,
            I => \N__46651\
        );

    \I__10937\ : CascadeMux
    port map (
            O => \N__46654\,
            I => \N__46648\
        );

    \I__10936\ : InMux
    port map (
            O => \N__46651\,
            I => \N__46643\
        );

    \I__10935\ : InMux
    port map (
            O => \N__46648\,
            I => \N__46643\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__46643\,
            I => \N__46639\
        );

    \I__10933\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46636\
        );

    \I__10932\ : Span4Mux_h
    port map (
            O => \N__46639\,
            I => \N__46633\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__46636\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__10930\ : Odrv4
    port map (
            O => \N__46633\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__10929\ : CascadeMux
    port map (
            O => \N__46628\,
            I => \N__46624\
        );

    \I__10928\ : CascadeMux
    port map (
            O => \N__46627\,
            I => \N__46621\
        );

    \I__10927\ : InMux
    port map (
            O => \N__46624\,
            I => \N__46617\
        );

    \I__10926\ : InMux
    port map (
            O => \N__46621\,
            I => \N__46612\
        );

    \I__10925\ : InMux
    port map (
            O => \N__46620\,
            I => \N__46612\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__46617\,
            I => \N__46609\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__46612\,
            I => \N__46606\
        );

    \I__10922\ : Span4Mux_h
    port map (
            O => \N__46609\,
            I => \N__46602\
        );

    \I__10921\ : Span4Mux_h
    port map (
            O => \N__46606\,
            I => \N__46599\
        );

    \I__10920\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46596\
        );

    \I__10919\ : Odrv4
    port map (
            O => \N__46602\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10918\ : Odrv4
    port map (
            O => \N__46599\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__46596\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10916\ : InMux
    port map (
            O => \N__46589\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__10915\ : InMux
    port map (
            O => \N__46586\,
            I => \N__46580\
        );

    \I__10914\ : InMux
    port map (
            O => \N__46585\,
            I => \N__46580\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__46580\,
            I => \N__46576\
        );

    \I__10912\ : InMux
    port map (
            O => \N__46579\,
            I => \N__46573\
        );

    \I__10911\ : Span4Mux_h
    port map (
            O => \N__46576\,
            I => \N__46570\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__46573\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__10909\ : Odrv4
    port map (
            O => \N__46570\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__10908\ : CascadeMux
    port map (
            O => \N__46565\,
            I => \N__46562\
        );

    \I__10907\ : InMux
    port map (
            O => \N__46562\,
            I => \N__46559\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__46559\,
            I => \N__46554\
        );

    \I__10905\ : InMux
    port map (
            O => \N__46558\,
            I => \N__46551\
        );

    \I__10904\ : InMux
    port map (
            O => \N__46557\,
            I => \N__46548\
        );

    \I__10903\ : Span4Mux_v
    port map (
            O => \N__46554\,
            I => \N__46543\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__46551\,
            I => \N__46543\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__46548\,
            I => \N__46539\
        );

    \I__10900\ : Span4Mux_h
    port map (
            O => \N__46543\,
            I => \N__46536\
        );

    \I__10899\ : InMux
    port map (
            O => \N__46542\,
            I => \N__46533\
        );

    \I__10898\ : Odrv12
    port map (
            O => \N__46539\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10897\ : Odrv4
    port map (
            O => \N__46536\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__46533\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10895\ : InMux
    port map (
            O => \N__46526\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__10894\ : CascadeMux
    port map (
            O => \N__46523\,
            I => \N__46520\
        );

    \I__10893\ : InMux
    port map (
            O => \N__46520\,
            I => \N__46516\
        );

    \I__10892\ : InMux
    port map (
            O => \N__46519\,
            I => \N__46513\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__46516\,
            I => \N__46509\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__46513\,
            I => \N__46506\
        );

    \I__10889\ : InMux
    port map (
            O => \N__46512\,
            I => \N__46503\
        );

    \I__10888\ : Span4Mux_h
    port map (
            O => \N__46509\,
            I => \N__46500\
        );

    \I__10887\ : Span4Mux_h
    port map (
            O => \N__46506\,
            I => \N__46497\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__46503\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__10885\ : Odrv4
    port map (
            O => \N__46500\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__10884\ : Odrv4
    port map (
            O => \N__46497\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__10883\ : CascadeMux
    port map (
            O => \N__46490\,
            I => \N__46487\
        );

    \I__10882\ : InMux
    port map (
            O => \N__46487\,
            I => \N__46484\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__46484\,
            I => \N__46479\
        );

    \I__10880\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46474\
        );

    \I__10879\ : InMux
    port map (
            O => \N__46482\,
            I => \N__46474\
        );

    \I__10878\ : Span4Mux_v
    port map (
            O => \N__46479\,
            I => \N__46468\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__46474\,
            I => \N__46468\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46465\
        );

    \I__10875\ : Odrv4
    port map (
            O => \N__46468\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__46465\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10873\ : InMux
    port map (
            O => \N__46460\,
            I => \bfn_18_20_0_\
        );

    \I__10872\ : CascadeMux
    port map (
            O => \N__46457\,
            I => \N__46454\
        );

    \I__10871\ : InMux
    port map (
            O => \N__46454\,
            I => \N__46450\
        );

    \I__10870\ : InMux
    port map (
            O => \N__46453\,
            I => \N__46447\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__46450\,
            I => \N__46443\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__46447\,
            I => \N__46440\
        );

    \I__10867\ : InMux
    port map (
            O => \N__46446\,
            I => \N__46437\
        );

    \I__10866\ : Span4Mux_h
    port map (
            O => \N__46443\,
            I => \N__46434\
        );

    \I__10865\ : Span4Mux_h
    port map (
            O => \N__46440\,
            I => \N__46431\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__46437\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10863\ : Odrv4
    port map (
            O => \N__46434\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10862\ : Odrv4
    port map (
            O => \N__46431\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10861\ : InMux
    port map (
            O => \N__46424\,
            I => \N__46420\
        );

    \I__10860\ : InMux
    port map (
            O => \N__46423\,
            I => \N__46416\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__46420\,
            I => \N__46413\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46419\,
            I => \N__46409\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__46416\,
            I => \N__46404\
        );

    \I__10856\ : Span12Mux_v
    port map (
            O => \N__46413\,
            I => \N__46404\
        );

    \I__10855\ : InMux
    port map (
            O => \N__46412\,
            I => \N__46401\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__46409\,
            I => \N__46398\
        );

    \I__10853\ : Odrv12
    port map (
            O => \N__46404\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__46401\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10851\ : Odrv4
    port map (
            O => \N__46398\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10850\ : InMux
    port map (
            O => \N__46391\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__10849\ : CascadeMux
    port map (
            O => \N__46388\,
            I => \N__46385\
        );

    \I__10848\ : InMux
    port map (
            O => \N__46385\,
            I => \N__46380\
        );

    \I__10847\ : InMux
    port map (
            O => \N__46384\,
            I => \N__46377\
        );

    \I__10846\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46374\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__46380\,
            I => \N__46369\
        );

    \I__10844\ : LocalMux
    port map (
            O => \N__46377\,
            I => \N__46369\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__46374\,
            I => \N__46364\
        );

    \I__10842\ : Span4Mux_v
    port map (
            O => \N__46369\,
            I => \N__46364\
        );

    \I__10841\ : Odrv4
    port map (
            O => \N__46364\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__10840\ : CascadeMux
    port map (
            O => \N__46361\,
            I => \N__46358\
        );

    \I__10839\ : InMux
    port map (
            O => \N__46358\,
            I => \N__46355\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__46355\,
            I => \N__46352\
        );

    \I__10837\ : Span4Mux_h
    port map (
            O => \N__46352\,
            I => \N__46348\
        );

    \I__10836\ : InMux
    port map (
            O => \N__46351\,
            I => \N__46345\
        );

    \I__10835\ : Span4Mux_h
    port map (
            O => \N__46348\,
            I => \N__46340\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__46345\,
            I => \N__46337\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46344\,
            I => \N__46334\
        );

    \I__10832\ : InMux
    port map (
            O => \N__46343\,
            I => \N__46331\
        );

    \I__10831\ : Odrv4
    port map (
            O => \N__46340\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10830\ : Odrv12
    port map (
            O => \N__46337\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__46334\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__46331\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__10827\ : InMux
    port map (
            O => \N__46322\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__10826\ : InMux
    port map (
            O => \N__46319\,
            I => \N__46313\
        );

    \I__10825\ : InMux
    port map (
            O => \N__46318\,
            I => \N__46313\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__46313\,
            I => \N__46309\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46312\,
            I => \N__46306\
        );

    \I__10822\ : Span4Mux_v
    port map (
            O => \N__46309\,
            I => \N__46303\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__46306\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__10820\ : Odrv4
    port map (
            O => \N__46303\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__10819\ : InMux
    port map (
            O => \N__46298\,
            I => \N__46295\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__46295\,
            I => \N__46289\
        );

    \I__10817\ : InMux
    port map (
            O => \N__46294\,
            I => \N__46284\
        );

    \I__10816\ : InMux
    port map (
            O => \N__46293\,
            I => \N__46284\
        );

    \I__10815\ : InMux
    port map (
            O => \N__46292\,
            I => \N__46281\
        );

    \I__10814\ : Span4Mux_v
    port map (
            O => \N__46289\,
            I => \N__46276\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__46284\,
            I => \N__46276\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__46281\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10811\ : Odrv4
    port map (
            O => \N__46276\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10810\ : InMux
    port map (
            O => \N__46271\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__10809\ : CascadeMux
    port map (
            O => \N__46268\,
            I => \N__46265\
        );

    \I__10808\ : InMux
    port map (
            O => \N__46265\,
            I => \N__46261\
        );

    \I__10807\ : InMux
    port map (
            O => \N__46264\,
            I => \N__46258\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__46261\,
            I => \N__46252\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46258\,
            I => \N__46252\
        );

    \I__10804\ : InMux
    port map (
            O => \N__46257\,
            I => \N__46249\
        );

    \I__10803\ : Span4Mux_h
    port map (
            O => \N__46252\,
            I => \N__46246\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__46249\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__10801\ : Odrv4
    port map (
            O => \N__46246\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__10800\ : CascadeMux
    port map (
            O => \N__46241\,
            I => \N__46238\
        );

    \I__10799\ : InMux
    port map (
            O => \N__46238\,
            I => \N__46235\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__46235\,
            I => \N__46231\
        );

    \I__10797\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46228\
        );

    \I__10796\ : Span4Mux_h
    port map (
            O => \N__46231\,
            I => \N__46222\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__46228\,
            I => \N__46222\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46227\,
            I => \N__46219\
        );

    \I__10793\ : Span4Mux_v
    port map (
            O => \N__46222\,
            I => \N__46216\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__46219\,
            I => \N__46212\
        );

    \I__10791\ : Span4Mux_h
    port map (
            O => \N__46216\,
            I => \N__46209\
        );

    \I__10790\ : InMux
    port map (
            O => \N__46215\,
            I => \N__46206\
        );

    \I__10789\ : Odrv12
    port map (
            O => \N__46212\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10788\ : Odrv4
    port map (
            O => \N__46209\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__46206\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10786\ : InMux
    port map (
            O => \N__46199\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__10785\ : CascadeMux
    port map (
            O => \N__46196\,
            I => \N__46192\
        );

    \I__10784\ : CascadeMux
    port map (
            O => \N__46195\,
            I => \N__46189\
        );

    \I__10783\ : InMux
    port map (
            O => \N__46192\,
            I => \N__46184\
        );

    \I__10782\ : InMux
    port map (
            O => \N__46189\,
            I => \N__46184\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46184\,
            I => \N__46180\
        );

    \I__10780\ : InMux
    port map (
            O => \N__46183\,
            I => \N__46177\
        );

    \I__10779\ : Span4Mux_h
    port map (
            O => \N__46180\,
            I => \N__46174\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__46177\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__10777\ : Odrv4
    port map (
            O => \N__46174\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__10776\ : CascadeMux
    port map (
            O => \N__46169\,
            I => \N__46166\
        );

    \I__10775\ : InMux
    port map (
            O => \N__46166\,
            I => \N__46161\
        );

    \I__10774\ : InMux
    port map (
            O => \N__46165\,
            I => \N__46158\
        );

    \I__10773\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46155\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__46161\,
            I => \N__46151\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__46158\,
            I => \N__46146\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46155\,
            I => \N__46146\
        );

    \I__10769\ : InMux
    port map (
            O => \N__46154\,
            I => \N__46143\
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__46151\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__10767\ : Odrv12
    port map (
            O => \N__46146\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__46143\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__10765\ : InMux
    port map (
            O => \N__46136\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__10764\ : InMux
    port map (
            O => \N__46133\,
            I => \N__46127\
        );

    \I__10763\ : InMux
    port map (
            O => \N__46132\,
            I => \N__46127\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__46127\,
            I => \N__46123\
        );

    \I__10761\ : InMux
    port map (
            O => \N__46126\,
            I => \N__46120\
        );

    \I__10760\ : Span4Mux_h
    port map (
            O => \N__46123\,
            I => \N__46117\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46120\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__10758\ : Odrv4
    port map (
            O => \N__46117\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__10757\ : CascadeMux
    port map (
            O => \N__46112\,
            I => \N__46107\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46111\,
            I => \N__46102\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46110\,
            I => \N__46102\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46107\,
            I => \N__46099\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__46102\,
            I => \N__46096\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__46099\,
            I => \N__46092\
        );

    \I__10751\ : Span4Mux_v
    port map (
            O => \N__46096\,
            I => \N__46089\
        );

    \I__10750\ : InMux
    port map (
            O => \N__46095\,
            I => \N__46086\
        );

    \I__10749\ : Odrv4
    port map (
            O => \N__46092\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10748\ : Odrv4
    port map (
            O => \N__46089\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10747\ : LocalMux
    port map (
            O => \N__46086\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46079\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46076\,
            I => \N__46070\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46075\,
            I => \N__46070\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__46070\,
            I => \N__46066\
        );

    \I__10742\ : InMux
    port map (
            O => \N__46069\,
            I => \N__46063\
        );

    \I__10741\ : Span4Mux_h
    port map (
            O => \N__46066\,
            I => \N__46060\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__46063\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__10739\ : Odrv4
    port map (
            O => \N__46060\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__10738\ : InMux
    port map (
            O => \N__46055\,
            I => \N__46051\
        );

    \I__10737\ : InMux
    port map (
            O => \N__46054\,
            I => \N__46047\
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__46051\,
            I => \N__46043\
        );

    \I__10735\ : InMux
    port map (
            O => \N__46050\,
            I => \N__46040\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__46047\,
            I => \N__46037\
        );

    \I__10733\ : InMux
    port map (
            O => \N__46046\,
            I => \N__46034\
        );

    \I__10732\ : Span4Mux_v
    port map (
            O => \N__46043\,
            I => \N__46029\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__46040\,
            I => \N__46029\
        );

    \I__10730\ : Odrv4
    port map (
            O => \N__46037\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__46034\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10728\ : Odrv4
    port map (
            O => \N__46029\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10727\ : InMux
    port map (
            O => \N__46022\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__10726\ : InMux
    port map (
            O => \N__46019\,
            I => \N__46015\
        );

    \I__10725\ : InMux
    port map (
            O => \N__46018\,
            I => \N__46012\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__46015\,
            I => \N__46009\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__46012\,
            I => \N__46005\
        );

    \I__10722\ : Span4Mux_v
    port map (
            O => \N__46009\,
            I => \N__46002\
        );

    \I__10721\ : InMux
    port map (
            O => \N__46008\,
            I => \N__45999\
        );

    \I__10720\ : Span4Mux_h
    port map (
            O => \N__46005\,
            I => \N__45996\
        );

    \I__10719\ : Odrv4
    port map (
            O => \N__46002\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__45999\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__10717\ : Odrv4
    port map (
            O => \N__45996\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__10716\ : CascadeMux
    port map (
            O => \N__45989\,
            I => \N__45986\
        );

    \I__10715\ : InMux
    port map (
            O => \N__45986\,
            I => \N__45979\
        );

    \I__10714\ : InMux
    port map (
            O => \N__45985\,
            I => \N__45979\
        );

    \I__10713\ : InMux
    port map (
            O => \N__45984\,
            I => \N__45976\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__45979\,
            I => \N__45972\
        );

    \I__10711\ : LocalMux
    port map (
            O => \N__45976\,
            I => \N__45969\
        );

    \I__10710\ : InMux
    port map (
            O => \N__45975\,
            I => \N__45966\
        );

    \I__10709\ : Span4Mux_v
    port map (
            O => \N__45972\,
            I => \N__45963\
        );

    \I__10708\ : Span4Mux_h
    port map (
            O => \N__45969\,
            I => \N__45960\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__45966\,
            I => \N__45957\
        );

    \I__10706\ : Odrv4
    port map (
            O => \N__45963\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10705\ : Odrv4
    port map (
            O => \N__45960\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10704\ : Odrv12
    port map (
            O => \N__45957\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10703\ : InMux
    port map (
            O => \N__45950\,
            I => \N__45947\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__45947\,
            I => \N__45943\
        );

    \I__10701\ : InMux
    port map (
            O => \N__45946\,
            I => \N__45940\
        );

    \I__10700\ : Span4Mux_v
    port map (
            O => \N__45943\,
            I => \N__45937\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__45940\,
            I => \N__45933\
        );

    \I__10698\ : Span4Mux_v
    port map (
            O => \N__45937\,
            I => \N__45930\
        );

    \I__10697\ : InMux
    port map (
            O => \N__45936\,
            I => \N__45927\
        );

    \I__10696\ : Span4Mux_h
    port map (
            O => \N__45933\,
            I => \N__45924\
        );

    \I__10695\ : Odrv4
    port map (
            O => \N__45930\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__45927\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10693\ : Odrv4
    port map (
            O => \N__45924\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10692\ : CascadeMux
    port map (
            O => \N__45917\,
            I => \N__45912\
        );

    \I__10691\ : InMux
    port map (
            O => \N__45916\,
            I => \N__45909\
        );

    \I__10690\ : InMux
    port map (
            O => \N__45915\,
            I => \N__45906\
        );

    \I__10689\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45903\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__45909\,
            I => \N__45900\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__45906\,
            I => \N__45894\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__45903\,
            I => \N__45894\
        );

    \I__10685\ : Span4Mux_h
    port map (
            O => \N__45900\,
            I => \N__45891\
        );

    \I__10684\ : InMux
    port map (
            O => \N__45899\,
            I => \N__45888\
        );

    \I__10683\ : Span12Mux_v
    port map (
            O => \N__45894\,
            I => \N__45885\
        );

    \I__10682\ : Span4Mux_h
    port map (
            O => \N__45891\,
            I => \N__45882\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__45888\,
            I => \N__45879\
        );

    \I__10680\ : Odrv12
    port map (
            O => \N__45885\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__10679\ : Odrv4
    port map (
            O => \N__45882\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__10678\ : Odrv12
    port map (
            O => \N__45879\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__10677\ : InMux
    port map (
            O => \N__45872\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__10676\ : CascadeMux
    port map (
            O => \N__45869\,
            I => \N__45865\
        );

    \I__10675\ : CascadeMux
    port map (
            O => \N__45868\,
            I => \N__45862\
        );

    \I__10674\ : InMux
    port map (
            O => \N__45865\,
            I => \N__45856\
        );

    \I__10673\ : InMux
    port map (
            O => \N__45862\,
            I => \N__45856\
        );

    \I__10672\ : InMux
    port map (
            O => \N__45861\,
            I => \N__45853\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__45856\,
            I => \N__45850\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__45853\,
            I => \N__45845\
        );

    \I__10669\ : Span4Mux_v
    port map (
            O => \N__45850\,
            I => \N__45845\
        );

    \I__10668\ : Odrv4
    port map (
            O => \N__45845\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__10667\ : InMux
    port map (
            O => \N__45842\,
            I => \N__45839\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__45839\,
            I => \N__45833\
        );

    \I__10665\ : InMux
    port map (
            O => \N__45838\,
            I => \N__45830\
        );

    \I__10664\ : InMux
    port map (
            O => \N__45837\,
            I => \N__45827\
        );

    \I__10663\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45824\
        );

    \I__10662\ : Span4Mux_h
    port map (
            O => \N__45833\,
            I => \N__45821\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__45830\,
            I => \N__45818\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__45827\,
            I => \N__45813\
        );

    \I__10659\ : LocalMux
    port map (
            O => \N__45824\,
            I => \N__45813\
        );

    \I__10658\ : Span4Mux_v
    port map (
            O => \N__45821\,
            I => \N__45810\
        );

    \I__10657\ : Span4Mux_h
    port map (
            O => \N__45818\,
            I => \N__45807\
        );

    \I__10656\ : Span4Mux_v
    port map (
            O => \N__45813\,
            I => \N__45804\
        );

    \I__10655\ : Odrv4
    port map (
            O => \N__45810\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__10654\ : Odrv4
    port map (
            O => \N__45807\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__10653\ : Odrv4
    port map (
            O => \N__45804\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__10652\ : InMux
    port map (
            O => \N__45797\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__10651\ : CascadeMux
    port map (
            O => \N__45794\,
            I => \N__45790\
        );

    \I__10650\ : CascadeMux
    port map (
            O => \N__45793\,
            I => \N__45787\
        );

    \I__10649\ : InMux
    port map (
            O => \N__45790\,
            I => \N__45782\
        );

    \I__10648\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45782\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__45782\,
            I => \N__45778\
        );

    \I__10646\ : InMux
    port map (
            O => \N__45781\,
            I => \N__45775\
        );

    \I__10645\ : Span4Mux_v
    port map (
            O => \N__45778\,
            I => \N__45772\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__45775\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__10643\ : Odrv4
    port map (
            O => \N__45772\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__10642\ : CascadeMux
    port map (
            O => \N__45767\,
            I => \N__45764\
        );

    \I__10641\ : InMux
    port map (
            O => \N__45764\,
            I => \N__45758\
        );

    \I__10640\ : InMux
    port map (
            O => \N__45763\,
            I => \N__45758\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__45758\,
            I => \N__45753\
        );

    \I__10638\ : InMux
    port map (
            O => \N__45757\,
            I => \N__45750\
        );

    \I__10637\ : InMux
    port map (
            O => \N__45756\,
            I => \N__45747\
        );

    \I__10636\ : Span4Mux_h
    port map (
            O => \N__45753\,
            I => \N__45744\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__45750\,
            I => \N__45741\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__45747\,
            I => \N__45738\
        );

    \I__10633\ : Span4Mux_v
    port map (
            O => \N__45744\,
            I => \N__45735\
        );

    \I__10632\ : Span4Mux_h
    port map (
            O => \N__45741\,
            I => \N__45732\
        );

    \I__10631\ : Span4Mux_v
    port map (
            O => \N__45738\,
            I => \N__45729\
        );

    \I__10630\ : Odrv4
    port map (
            O => \N__45735\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__10629\ : Odrv4
    port map (
            O => \N__45732\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__10628\ : Odrv4
    port map (
            O => \N__45729\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__10627\ : InMux
    port map (
            O => \N__45722\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__10626\ : CascadeMux
    port map (
            O => \N__45719\,
            I => \N__45716\
        );

    \I__10625\ : InMux
    port map (
            O => \N__45716\,
            I => \N__45712\
        );

    \I__10624\ : InMux
    port map (
            O => \N__45715\,
            I => \N__45709\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__45712\,
            I => \N__45703\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__45709\,
            I => \N__45703\
        );

    \I__10621\ : InMux
    port map (
            O => \N__45708\,
            I => \N__45700\
        );

    \I__10620\ : Span4Mux_h
    port map (
            O => \N__45703\,
            I => \N__45697\
        );

    \I__10619\ : LocalMux
    port map (
            O => \N__45700\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__10618\ : Odrv4
    port map (
            O => \N__45697\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__10617\ : CascadeMux
    port map (
            O => \N__45692\,
            I => \N__45688\
        );

    \I__10616\ : InMux
    port map (
            O => \N__45691\,
            I => \N__45683\
        );

    \I__10615\ : InMux
    port map (
            O => \N__45688\,
            I => \N__45683\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__45683\,
            I => \N__45679\
        );

    \I__10613\ : InMux
    port map (
            O => \N__45682\,
            I => \N__45676\
        );

    \I__10612\ : Span4Mux_h
    port map (
            O => \N__45679\,
            I => \N__45673\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__45676\,
            I => \N__45670\
        );

    \I__10610\ : Span4Mux_v
    port map (
            O => \N__45673\,
            I => \N__45666\
        );

    \I__10609\ : Span4Mux_h
    port map (
            O => \N__45670\,
            I => \N__45663\
        );

    \I__10608\ : InMux
    port map (
            O => \N__45669\,
            I => \N__45660\
        );

    \I__10607\ : Odrv4
    port map (
            O => \N__45666\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10606\ : Odrv4
    port map (
            O => \N__45663\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__45660\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10604\ : InMux
    port map (
            O => \N__45653\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__10603\ : CascadeMux
    port map (
            O => \N__45650\,
            I => \N__45647\
        );

    \I__10602\ : InMux
    port map (
            O => \N__45647\,
            I => \N__45643\
        );

    \I__10601\ : InMux
    port map (
            O => \N__45646\,
            I => \N__45640\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__45643\,
            I => \N__45634\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__45640\,
            I => \N__45634\
        );

    \I__10598\ : InMux
    port map (
            O => \N__45639\,
            I => \N__45631\
        );

    \I__10597\ : Span4Mux_h
    port map (
            O => \N__45634\,
            I => \N__45628\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__45631\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__10595\ : Odrv4
    port map (
            O => \N__45628\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__10594\ : CascadeMux
    port map (
            O => \N__45623\,
            I => \N__45619\
        );

    \I__10593\ : CascadeMux
    port map (
            O => \N__45622\,
            I => \N__45616\
        );

    \I__10592\ : InMux
    port map (
            O => \N__45619\,
            I => \N__45611\
        );

    \I__10591\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45611\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__45611\,
            I => \N__45607\
        );

    \I__10589\ : InMux
    port map (
            O => \N__45610\,
            I => \N__45604\
        );

    \I__10588\ : Span4Mux_h
    port map (
            O => \N__45607\,
            I => \N__45600\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__45604\,
            I => \N__45597\
        );

    \I__10586\ : InMux
    port map (
            O => \N__45603\,
            I => \N__45594\
        );

    \I__10585\ : Span4Mux_v
    port map (
            O => \N__45600\,
            I => \N__45591\
        );

    \I__10584\ : Span4Mux_h
    port map (
            O => \N__45597\,
            I => \N__45588\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__45594\,
            I => \N__45585\
        );

    \I__10582\ : Odrv4
    port map (
            O => \N__45591\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__10581\ : Odrv4
    port map (
            O => \N__45588\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__10580\ : Odrv12
    port map (
            O => \N__45585\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__10579\ : InMux
    port map (
            O => \N__45578\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__10578\ : CascadeMux
    port map (
            O => \N__45575\,
            I => \N__45572\
        );

    \I__10577\ : InMux
    port map (
            O => \N__45572\,
            I => \N__45568\
        );

    \I__10576\ : InMux
    port map (
            O => \N__45571\,
            I => \N__45565\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__45568\,
            I => \N__45559\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__45565\,
            I => \N__45559\
        );

    \I__10573\ : InMux
    port map (
            O => \N__45564\,
            I => \N__45556\
        );

    \I__10572\ : Span4Mux_h
    port map (
            O => \N__45559\,
            I => \N__45553\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__45556\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__10570\ : Odrv4
    port map (
            O => \N__45553\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__10569\ : CascadeMux
    port map (
            O => \N__45548\,
            I => \N__45545\
        );

    \I__10568\ : InMux
    port map (
            O => \N__45545\,
            I => \N__45540\
        );

    \I__10567\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45535\
        );

    \I__10566\ : InMux
    port map (
            O => \N__45543\,
            I => \N__45535\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__45540\,
            I => \N__45530\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__45535\,
            I => \N__45530\
        );

    \I__10563\ : Span12Mux_v
    port map (
            O => \N__45530\,
            I => \N__45526\
        );

    \I__10562\ : InMux
    port map (
            O => \N__45529\,
            I => \N__45523\
        );

    \I__10561\ : Odrv12
    port map (
            O => \N__45526\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__45523\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10559\ : InMux
    port map (
            O => \N__45518\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__10558\ : CascadeMux
    port map (
            O => \N__45515\,
            I => \N__45512\
        );

    \I__10557\ : InMux
    port map (
            O => \N__45512\,
            I => \N__45508\
        );

    \I__10556\ : InMux
    port map (
            O => \N__45511\,
            I => \N__45505\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__45508\,
            I => \N__45499\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__45505\,
            I => \N__45499\
        );

    \I__10553\ : InMux
    port map (
            O => \N__45504\,
            I => \N__45496\
        );

    \I__10552\ : Span4Mux_h
    port map (
            O => \N__45499\,
            I => \N__45493\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__45496\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__10550\ : Odrv4
    port map (
            O => \N__45493\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__10549\ : CascadeMux
    port map (
            O => \N__45488\,
            I => \N__45485\
        );

    \I__10548\ : InMux
    port map (
            O => \N__45485\,
            I => \N__45482\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__45482\,
            I => \N__45479\
        );

    \I__10546\ : Span4Mux_h
    port map (
            O => \N__45479\,
            I => \N__45474\
        );

    \I__10545\ : InMux
    port map (
            O => \N__45478\,
            I => \N__45471\
        );

    \I__10544\ : InMux
    port map (
            O => \N__45477\,
            I => \N__45467\
        );

    \I__10543\ : Span4Mux_h
    port map (
            O => \N__45474\,
            I => \N__45464\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__45471\,
            I => \N__45461\
        );

    \I__10541\ : InMux
    port map (
            O => \N__45470\,
            I => \N__45458\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__45467\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10539\ : Odrv4
    port map (
            O => \N__45464\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10538\ : Odrv12
    port map (
            O => \N__45461\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__45458\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10536\ : InMux
    port map (
            O => \N__45449\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__10535\ : CascadeMux
    port map (
            O => \N__45446\,
            I => \N__45443\
        );

    \I__10534\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45440\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__45440\,
            I => \N__45437\
        );

    \I__10532\ : Span4Mux_h
    port map (
            O => \N__45437\,
            I => \N__45434\
        );

    \I__10531\ : Span4Mux_v
    port map (
            O => \N__45434\,
            I => \N__45431\
        );

    \I__10530\ : Odrv4
    port map (
            O => \N__45431\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__10529\ : CascadeMux
    port map (
            O => \N__45428\,
            I => \N__45425\
        );

    \I__10528\ : InMux
    port map (
            O => \N__45425\,
            I => \N__45421\
        );

    \I__10527\ : CascadeMux
    port map (
            O => \N__45424\,
            I => \N__45418\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__45421\,
            I => \N__45414\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45418\,
            I => \N__45411\
        );

    \I__10524\ : InMux
    port map (
            O => \N__45417\,
            I => \N__45408\
        );

    \I__10523\ : Odrv4
    port map (
            O => \N__45414\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__45411\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__45408\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10520\ : CascadeMux
    port map (
            O => \N__45401\,
            I => \N__45398\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45398\,
            I => \N__45395\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__45395\,
            I => \N__45392\
        );

    \I__10517\ : Span4Mux_v
    port map (
            O => \N__45392\,
            I => \N__45389\
        );

    \I__10516\ : Span4Mux_h
    port map (
            O => \N__45389\,
            I => \N__45386\
        );

    \I__10515\ : Odrv4
    port map (
            O => \N__45386\,
            I => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\
        );

    \I__10514\ : InMux
    port map (
            O => \N__45383\,
            I => \N__45380\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__45380\,
            I => \N__45377\
        );

    \I__10512\ : Odrv4
    port map (
            O => \N__45377\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__10511\ : InMux
    port map (
            O => \N__45374\,
            I => \N__45371\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__45371\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__10509\ : InMux
    port map (
            O => \N__45368\,
            I => \N__45363\
        );

    \I__10508\ : InMux
    port map (
            O => \N__45367\,
            I => \N__45360\
        );

    \I__10507\ : InMux
    port map (
            O => \N__45366\,
            I => \N__45357\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__45363\,
            I => \N__45354\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__45360\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__45357\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__10503\ : Odrv4
    port map (
            O => \N__45354\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__10502\ : CascadeMux
    port map (
            O => \N__45347\,
            I => \N__45344\
        );

    \I__10501\ : InMux
    port map (
            O => \N__45344\,
            I => \N__45341\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__45341\,
            I => \N__45338\
        );

    \I__10499\ : Span4Mux_v
    port map (
            O => \N__45338\,
            I => \N__45335\
        );

    \I__10498\ : Span4Mux_h
    port map (
            O => \N__45335\,
            I => \N__45332\
        );

    \I__10497\ : Odrv4
    port map (
            O => \N__45332\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__10496\ : InMux
    port map (
            O => \N__45329\,
            I => \N__45326\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__45326\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__10494\ : InMux
    port map (
            O => \N__45323\,
            I => \N__45320\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__45320\,
            I => \N__45317\
        );

    \I__10492\ : Span4Mux_v
    port map (
            O => \N__45317\,
            I => \N__45312\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45316\,
            I => \N__45309\
        );

    \I__10490\ : InMux
    port map (
            O => \N__45315\,
            I => \N__45306\
        );

    \I__10489\ : Span4Mux_h
    port map (
            O => \N__45312\,
            I => \N__45303\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__45309\,
            I => \N__45300\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__45306\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__10486\ : Odrv4
    port map (
            O => \N__45303\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__10485\ : Odrv4
    port map (
            O => \N__45300\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__10484\ : CascadeMux
    port map (
            O => \N__45293\,
            I => \N__45284\
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__45292\,
            I => \N__45281\
        );

    \I__10482\ : CascadeMux
    port map (
            O => \N__45291\,
            I => \N__45275\
        );

    \I__10481\ : CascadeMux
    port map (
            O => \N__45290\,
            I => \N__45272\
        );

    \I__10480\ : CascadeMux
    port map (
            O => \N__45289\,
            I => \N__45268\
        );

    \I__10479\ : CascadeMux
    port map (
            O => \N__45288\,
            I => \N__45260\
        );

    \I__10478\ : CascadeMux
    port map (
            O => \N__45287\,
            I => \N__45254\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45284\,
            I => \N__45248\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45281\,
            I => \N__45248\
        );

    \I__10475\ : CascadeMux
    port map (
            O => \N__45280\,
            I => \N__45245\
        );

    \I__10474\ : CascadeMux
    port map (
            O => \N__45279\,
            I => \N__45242\
        );

    \I__10473\ : CascadeMux
    port map (
            O => \N__45278\,
            I => \N__45238\
        );

    \I__10472\ : InMux
    port map (
            O => \N__45275\,
            I => \N__45227\
        );

    \I__10471\ : InMux
    port map (
            O => \N__45272\,
            I => \N__45227\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45271\,
            I => \N__45216\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45268\,
            I => \N__45216\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45267\,
            I => \N__45216\
        );

    \I__10467\ : InMux
    port map (
            O => \N__45266\,
            I => \N__45216\
        );

    \I__10466\ : InMux
    port map (
            O => \N__45265\,
            I => \N__45216\
        );

    \I__10465\ : CascadeMux
    port map (
            O => \N__45264\,
            I => \N__45212\
        );

    \I__10464\ : CascadeMux
    port map (
            O => \N__45263\,
            I => \N__45203\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45260\,
            I => \N__45195\
        );

    \I__10462\ : InMux
    port map (
            O => \N__45259\,
            I => \N__45190\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45258\,
            I => \N__45190\
        );

    \I__10460\ : InMux
    port map (
            O => \N__45257\,
            I => \N__45185\
        );

    \I__10459\ : InMux
    port map (
            O => \N__45254\,
            I => \N__45185\
        );

    \I__10458\ : CascadeMux
    port map (
            O => \N__45253\,
            I => \N__45182\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__45248\,
            I => \N__45173\
        );

    \I__10456\ : InMux
    port map (
            O => \N__45245\,
            I => \N__45170\
        );

    \I__10455\ : InMux
    port map (
            O => \N__45242\,
            I => \N__45163\
        );

    \I__10454\ : InMux
    port map (
            O => \N__45241\,
            I => \N__45163\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45238\,
            I => \N__45163\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45237\,
            I => \N__45152\
        );

    \I__10451\ : InMux
    port map (
            O => \N__45236\,
            I => \N__45152\
        );

    \I__10450\ : InMux
    port map (
            O => \N__45235\,
            I => \N__45152\
        );

    \I__10449\ : InMux
    port map (
            O => \N__45234\,
            I => \N__45152\
        );

    \I__10448\ : InMux
    port map (
            O => \N__45233\,
            I => \N__45152\
        );

    \I__10447\ : CascadeMux
    port map (
            O => \N__45232\,
            I => \N__45149\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45227\,
            I => \N__45120\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__45216\,
            I => \N__45120\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45215\,
            I => \N__45113\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45212\,
            I => \N__45113\
        );

    \I__10442\ : InMux
    port map (
            O => \N__45211\,
            I => \N__45113\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45210\,
            I => \N__45102\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45209\,
            I => \N__45102\
        );

    \I__10439\ : InMux
    port map (
            O => \N__45208\,
            I => \N__45102\
        );

    \I__10438\ : InMux
    port map (
            O => \N__45207\,
            I => \N__45102\
        );

    \I__10437\ : InMux
    port map (
            O => \N__45206\,
            I => \N__45102\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45203\,
            I => \N__45099\
        );

    \I__10435\ : CascadeMux
    port map (
            O => \N__45202\,
            I => \N__45095\
        );

    \I__10434\ : CascadeMux
    port map (
            O => \N__45201\,
            I => \N__45092\
        );

    \I__10433\ : InMux
    port map (
            O => \N__45200\,
            I => \N__45085\
        );

    \I__10432\ : InMux
    port map (
            O => \N__45199\,
            I => \N__45085\
        );

    \I__10431\ : InMux
    port map (
            O => \N__45198\,
            I => \N__45085\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__45195\,
            I => \N__45080\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__45190\,
            I => \N__45080\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45185\,
            I => \N__45077\
        );

    \I__10427\ : InMux
    port map (
            O => \N__45182\,
            I => \N__45074\
        );

    \I__10426\ : InMux
    port map (
            O => \N__45181\,
            I => \N__45071\
        );

    \I__10425\ : CascadeMux
    port map (
            O => \N__45180\,
            I => \N__45067\
        );

    \I__10424\ : CascadeMux
    port map (
            O => \N__45179\,
            I => \N__45062\
        );

    \I__10423\ : CascadeMux
    port map (
            O => \N__45178\,
            I => \N__45055\
        );

    \I__10422\ : CascadeMux
    port map (
            O => \N__45177\,
            I => \N__45052\
        );

    \I__10421\ : CascadeMux
    port map (
            O => \N__45176\,
            I => \N__45048\
        );

    \I__10420\ : Span4Mux_v
    port map (
            O => \N__45173\,
            I => \N__45032\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__45170\,
            I => \N__45032\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__45163\,
            I => \N__45032\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__45152\,
            I => \N__45032\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45149\,
            I => \N__45023\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45148\,
            I => \N__45023\
        );

    \I__10414\ : InMux
    port map (
            O => \N__45147\,
            I => \N__45023\
        );

    \I__10413\ : InMux
    port map (
            O => \N__45146\,
            I => \N__45023\
        );

    \I__10412\ : CascadeMux
    port map (
            O => \N__45145\,
            I => \N__45019\
        );

    \I__10411\ : CascadeMux
    port map (
            O => \N__45144\,
            I => \N__45015\
        );

    \I__10410\ : CascadeMux
    port map (
            O => \N__45143\,
            I => \N__45011\
        );

    \I__10409\ : CascadeMux
    port map (
            O => \N__45142\,
            I => \N__45005\
        );

    \I__10408\ : CascadeMux
    port map (
            O => \N__45141\,
            I => \N__45001\
        );

    \I__10407\ : CascadeMux
    port map (
            O => \N__45140\,
            I => \N__44997\
        );

    \I__10406\ : CascadeMux
    port map (
            O => \N__45139\,
            I => \N__44992\
        );

    \I__10405\ : CascadeMux
    port map (
            O => \N__45138\,
            I => \N__44988\
        );

    \I__10404\ : CascadeMux
    port map (
            O => \N__45137\,
            I => \N__44984\
        );

    \I__10403\ : CascadeMux
    port map (
            O => \N__45136\,
            I => \N__44980\
        );

    \I__10402\ : CascadeMux
    port map (
            O => \N__45135\,
            I => \N__44977\
        );

    \I__10401\ : CascadeMux
    port map (
            O => \N__45134\,
            I => \N__44973\
        );

    \I__10400\ : CascadeMux
    port map (
            O => \N__45133\,
            I => \N__44969\
        );

    \I__10399\ : CascadeMux
    port map (
            O => \N__45132\,
            I => \N__44965\
        );

    \I__10398\ : CascadeMux
    port map (
            O => \N__45131\,
            I => \N__44961\
        );

    \I__10397\ : CascadeMux
    port map (
            O => \N__45130\,
            I => \N__44957\
        );

    \I__10396\ : CascadeMux
    port map (
            O => \N__45129\,
            I => \N__44953\
        );

    \I__10395\ : CascadeMux
    port map (
            O => \N__45128\,
            I => \N__44949\
        );

    \I__10394\ : CascadeMux
    port map (
            O => \N__45127\,
            I => \N__44945\
        );

    \I__10393\ : CascadeMux
    port map (
            O => \N__45126\,
            I => \N__44941\
        );

    \I__10392\ : CascadeMux
    port map (
            O => \N__45125\,
            I => \N__44937\
        );

    \I__10391\ : Span4Mux_v
    port map (
            O => \N__45120\,
            I => \N__44931\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__45113\,
            I => \N__44931\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__45102\,
            I => \N__44928\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__45099\,
            I => \N__44925\
        );

    \I__10387\ : InMux
    port map (
            O => \N__45098\,
            I => \N__44922\
        );

    \I__10386\ : InMux
    port map (
            O => \N__45095\,
            I => \N__44917\
        );

    \I__10385\ : InMux
    port map (
            O => \N__45092\,
            I => \N__44917\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__45085\,
            I => \N__44914\
        );

    \I__10383\ : Span4Mux_v
    port map (
            O => \N__45080\,
            I => \N__44905\
        );

    \I__10382\ : Span4Mux_v
    port map (
            O => \N__45077\,
            I => \N__44905\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__45074\,
            I => \N__44905\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__45071\,
            I => \N__44905\
        );

    \I__10379\ : CascadeMux
    port map (
            O => \N__45070\,
            I => \N__44902\
        );

    \I__10378\ : InMux
    port map (
            O => \N__45067\,
            I => \N__44893\
        );

    \I__10377\ : InMux
    port map (
            O => \N__45066\,
            I => \N__44893\
        );

    \I__10376\ : InMux
    port map (
            O => \N__45065\,
            I => \N__44893\
        );

    \I__10375\ : InMux
    port map (
            O => \N__45062\,
            I => \N__44893\
        );

    \I__10374\ : InMux
    port map (
            O => \N__45061\,
            I => \N__44876\
        );

    \I__10373\ : InMux
    port map (
            O => \N__45060\,
            I => \N__44876\
        );

    \I__10372\ : InMux
    port map (
            O => \N__45059\,
            I => \N__44876\
        );

    \I__10371\ : InMux
    port map (
            O => \N__45058\,
            I => \N__44876\
        );

    \I__10370\ : InMux
    port map (
            O => \N__45055\,
            I => \N__44876\
        );

    \I__10369\ : InMux
    port map (
            O => \N__45052\,
            I => \N__44876\
        );

    \I__10368\ : InMux
    port map (
            O => \N__45051\,
            I => \N__44876\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45048\,
            I => \N__44876\
        );

    \I__10366\ : CascadeMux
    port map (
            O => \N__45047\,
            I => \N__44872\
        );

    \I__10365\ : CascadeMux
    port map (
            O => \N__45046\,
            I => \N__44868\
        );

    \I__10364\ : CascadeMux
    port map (
            O => \N__45045\,
            I => \N__44864\
        );

    \I__10363\ : CascadeMux
    port map (
            O => \N__45044\,
            I => \N__44860\
        );

    \I__10362\ : CascadeMux
    port map (
            O => \N__45043\,
            I => \N__44857\
        );

    \I__10361\ : CascadeMux
    port map (
            O => \N__45042\,
            I => \N__44853\
        );

    \I__10360\ : CascadeMux
    port map (
            O => \N__45041\,
            I => \N__44849\
        );

    \I__10359\ : Span4Mux_v
    port map (
            O => \N__45032\,
            I => \N__44843\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__45023\,
            I => \N__44843\
        );

    \I__10357\ : InMux
    port map (
            O => \N__45022\,
            I => \N__44828\
        );

    \I__10356\ : InMux
    port map (
            O => \N__45019\,
            I => \N__44828\
        );

    \I__10355\ : InMux
    port map (
            O => \N__45018\,
            I => \N__44828\
        );

    \I__10354\ : InMux
    port map (
            O => \N__45015\,
            I => \N__44828\
        );

    \I__10353\ : InMux
    port map (
            O => \N__45014\,
            I => \N__44828\
        );

    \I__10352\ : InMux
    port map (
            O => \N__45011\,
            I => \N__44828\
        );

    \I__10351\ : InMux
    port map (
            O => \N__45010\,
            I => \N__44828\
        );

    \I__10350\ : InMux
    port map (
            O => \N__45009\,
            I => \N__44811\
        );

    \I__10349\ : InMux
    port map (
            O => \N__45008\,
            I => \N__44811\
        );

    \I__10348\ : InMux
    port map (
            O => \N__45005\,
            I => \N__44811\
        );

    \I__10347\ : InMux
    port map (
            O => \N__45004\,
            I => \N__44811\
        );

    \I__10346\ : InMux
    port map (
            O => \N__45001\,
            I => \N__44811\
        );

    \I__10345\ : InMux
    port map (
            O => \N__45000\,
            I => \N__44811\
        );

    \I__10344\ : InMux
    port map (
            O => \N__44997\,
            I => \N__44811\
        );

    \I__10343\ : InMux
    port map (
            O => \N__44996\,
            I => \N__44811\
        );

    \I__10342\ : InMux
    port map (
            O => \N__44995\,
            I => \N__44794\
        );

    \I__10341\ : InMux
    port map (
            O => \N__44992\,
            I => \N__44794\
        );

    \I__10340\ : InMux
    port map (
            O => \N__44991\,
            I => \N__44794\
        );

    \I__10339\ : InMux
    port map (
            O => \N__44988\,
            I => \N__44794\
        );

    \I__10338\ : InMux
    port map (
            O => \N__44987\,
            I => \N__44794\
        );

    \I__10337\ : InMux
    port map (
            O => \N__44984\,
            I => \N__44794\
        );

    \I__10336\ : InMux
    port map (
            O => \N__44983\,
            I => \N__44794\
        );

    \I__10335\ : InMux
    port map (
            O => \N__44980\,
            I => \N__44794\
        );

    \I__10334\ : InMux
    port map (
            O => \N__44977\,
            I => \N__44777\
        );

    \I__10333\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44777\
        );

    \I__10332\ : InMux
    port map (
            O => \N__44973\,
            I => \N__44777\
        );

    \I__10331\ : InMux
    port map (
            O => \N__44972\,
            I => \N__44777\
        );

    \I__10330\ : InMux
    port map (
            O => \N__44969\,
            I => \N__44777\
        );

    \I__10329\ : InMux
    port map (
            O => \N__44968\,
            I => \N__44777\
        );

    \I__10328\ : InMux
    port map (
            O => \N__44965\,
            I => \N__44777\
        );

    \I__10327\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44777\
        );

    \I__10326\ : InMux
    port map (
            O => \N__44961\,
            I => \N__44760\
        );

    \I__10325\ : InMux
    port map (
            O => \N__44960\,
            I => \N__44760\
        );

    \I__10324\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44760\
        );

    \I__10323\ : InMux
    port map (
            O => \N__44956\,
            I => \N__44760\
        );

    \I__10322\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44760\
        );

    \I__10321\ : InMux
    port map (
            O => \N__44952\,
            I => \N__44760\
        );

    \I__10320\ : InMux
    port map (
            O => \N__44949\,
            I => \N__44760\
        );

    \I__10319\ : InMux
    port map (
            O => \N__44948\,
            I => \N__44760\
        );

    \I__10318\ : InMux
    port map (
            O => \N__44945\,
            I => \N__44747\
        );

    \I__10317\ : InMux
    port map (
            O => \N__44944\,
            I => \N__44747\
        );

    \I__10316\ : InMux
    port map (
            O => \N__44941\,
            I => \N__44747\
        );

    \I__10315\ : InMux
    port map (
            O => \N__44940\,
            I => \N__44747\
        );

    \I__10314\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44747\
        );

    \I__10313\ : InMux
    port map (
            O => \N__44936\,
            I => \N__44747\
        );

    \I__10312\ : Span4Mux_h
    port map (
            O => \N__44931\,
            I => \N__44744\
        );

    \I__10311\ : Span4Mux_v
    port map (
            O => \N__44928\,
            I => \N__44735\
        );

    \I__10310\ : Span4Mux_v
    port map (
            O => \N__44925\,
            I => \N__44735\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__44922\,
            I => \N__44735\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__44917\,
            I => \N__44735\
        );

    \I__10307\ : Span4Mux_v
    port map (
            O => \N__44914\,
            I => \N__44730\
        );

    \I__10306\ : Span4Mux_v
    port map (
            O => \N__44905\,
            I => \N__44730\
        );

    \I__10305\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44727\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__44893\,
            I => \N__44722\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__44876\,
            I => \N__44722\
        );

    \I__10302\ : InMux
    port map (
            O => \N__44875\,
            I => \N__44705\
        );

    \I__10301\ : InMux
    port map (
            O => \N__44872\,
            I => \N__44705\
        );

    \I__10300\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44705\
        );

    \I__10299\ : InMux
    port map (
            O => \N__44868\,
            I => \N__44705\
        );

    \I__10298\ : InMux
    port map (
            O => \N__44867\,
            I => \N__44705\
        );

    \I__10297\ : InMux
    port map (
            O => \N__44864\,
            I => \N__44705\
        );

    \I__10296\ : InMux
    port map (
            O => \N__44863\,
            I => \N__44705\
        );

    \I__10295\ : InMux
    port map (
            O => \N__44860\,
            I => \N__44705\
        );

    \I__10294\ : InMux
    port map (
            O => \N__44857\,
            I => \N__44692\
        );

    \I__10293\ : InMux
    port map (
            O => \N__44856\,
            I => \N__44692\
        );

    \I__10292\ : InMux
    port map (
            O => \N__44853\,
            I => \N__44692\
        );

    \I__10291\ : InMux
    port map (
            O => \N__44852\,
            I => \N__44692\
        );

    \I__10290\ : InMux
    port map (
            O => \N__44849\,
            I => \N__44692\
        );

    \I__10289\ : InMux
    port map (
            O => \N__44848\,
            I => \N__44692\
        );

    \I__10288\ : Sp12to4
    port map (
            O => \N__44843\,
            I => \N__44677\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__44828\,
            I => \N__44677\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__44811\,
            I => \N__44677\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__44794\,
            I => \N__44677\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__44777\,
            I => \N__44677\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__44760\,
            I => \N__44677\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__44747\,
            I => \N__44677\
        );

    \I__10281\ : Odrv4
    port map (
            O => \N__44744\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10280\ : Odrv4
    port map (
            O => \N__44735\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10279\ : Odrv4
    port map (
            O => \N__44730\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__44727\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10277\ : Odrv12
    port map (
            O => \N__44722\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__44705\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__44692\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10274\ : Odrv12
    port map (
            O => \N__44677\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10273\ : InMux
    port map (
            O => \N__44660\,
            I => \N__44639\
        );

    \I__10272\ : InMux
    port map (
            O => \N__44659\,
            I => \N__44639\
        );

    \I__10271\ : InMux
    port map (
            O => \N__44658\,
            I => \N__44630\
        );

    \I__10270\ : InMux
    port map (
            O => \N__44657\,
            I => \N__44630\
        );

    \I__10269\ : InMux
    port map (
            O => \N__44656\,
            I => \N__44630\
        );

    \I__10268\ : InMux
    port map (
            O => \N__44655\,
            I => \N__44630\
        );

    \I__10267\ : InMux
    port map (
            O => \N__44654\,
            I => \N__44615\
        );

    \I__10266\ : InMux
    port map (
            O => \N__44653\,
            I => \N__44612\
        );

    \I__10265\ : InMux
    port map (
            O => \N__44652\,
            I => \N__44606\
        );

    \I__10264\ : InMux
    port map (
            O => \N__44651\,
            I => \N__44595\
        );

    \I__10263\ : InMux
    port map (
            O => \N__44650\,
            I => \N__44595\
        );

    \I__10262\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44595\
        );

    \I__10261\ : InMux
    port map (
            O => \N__44648\,
            I => \N__44595\
        );

    \I__10260\ : InMux
    port map (
            O => \N__44647\,
            I => \N__44595\
        );

    \I__10259\ : InMux
    port map (
            O => \N__44646\,
            I => \N__44587\
        );

    \I__10258\ : InMux
    port map (
            O => \N__44645\,
            I => \N__44583\
        );

    \I__10257\ : InMux
    port map (
            O => \N__44644\,
            I => \N__44580\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__44639\,
            I => \N__44568\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__44630\,
            I => \N__44568\
        );

    \I__10254\ : InMux
    port map (
            O => \N__44629\,
            I => \N__44557\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44628\,
            I => \N__44557\
        );

    \I__10252\ : InMux
    port map (
            O => \N__44627\,
            I => \N__44557\
        );

    \I__10251\ : InMux
    port map (
            O => \N__44626\,
            I => \N__44557\
        );

    \I__10250\ : InMux
    port map (
            O => \N__44625\,
            I => \N__44557\
        );

    \I__10249\ : InMux
    port map (
            O => \N__44624\,
            I => \N__44554\
        );

    \I__10248\ : InMux
    port map (
            O => \N__44623\,
            I => \N__44547\
        );

    \I__10247\ : InMux
    port map (
            O => \N__44622\,
            I => \N__44547\
        );

    \I__10246\ : InMux
    port map (
            O => \N__44621\,
            I => \N__44547\
        );

    \I__10245\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44540\
        );

    \I__10244\ : InMux
    port map (
            O => \N__44619\,
            I => \N__44540\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44618\,
            I => \N__44540\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__44615\,
            I => \N__44535\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__44612\,
            I => \N__44535\
        );

    \I__10240\ : InMux
    port map (
            O => \N__44611\,
            I => \N__44531\
        );

    \I__10239\ : InMux
    port map (
            O => \N__44610\,
            I => \N__44528\
        );

    \I__10238\ : InMux
    port map (
            O => \N__44609\,
            I => \N__44525\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__44606\,
            I => \N__44520\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__44595\,
            I => \N__44520\
        );

    \I__10235\ : InMux
    port map (
            O => \N__44594\,
            I => \N__44509\
        );

    \I__10234\ : InMux
    port map (
            O => \N__44593\,
            I => \N__44509\
        );

    \I__10233\ : InMux
    port map (
            O => \N__44592\,
            I => \N__44509\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44591\,
            I => \N__44509\
        );

    \I__10231\ : InMux
    port map (
            O => \N__44590\,
            I => \N__44509\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__44587\,
            I => \N__44506\
        );

    \I__10229\ : InMux
    port map (
            O => \N__44586\,
            I => \N__44503\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__44583\,
            I => \N__44500\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__44580\,
            I => \N__44497\
        );

    \I__10226\ : InMux
    port map (
            O => \N__44579\,
            I => \N__44492\
        );

    \I__10225\ : InMux
    port map (
            O => \N__44578\,
            I => \N__44492\
        );

    \I__10224\ : InMux
    port map (
            O => \N__44577\,
            I => \N__44481\
        );

    \I__10223\ : InMux
    port map (
            O => \N__44576\,
            I => \N__44481\
        );

    \I__10222\ : InMux
    port map (
            O => \N__44575\,
            I => \N__44481\
        );

    \I__10221\ : InMux
    port map (
            O => \N__44574\,
            I => \N__44481\
        );

    \I__10220\ : InMux
    port map (
            O => \N__44573\,
            I => \N__44481\
        );

    \I__10219\ : Span4Mux_v
    port map (
            O => \N__44568\,
            I => \N__44471\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__44557\,
            I => \N__44471\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__44554\,
            I => \N__44466\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__44547\,
            I => \N__44466\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__44540\,
            I => \N__44458\
        );

    \I__10214\ : Span4Mux_v
    port map (
            O => \N__44535\,
            I => \N__44458\
        );

    \I__10213\ : InMux
    port map (
            O => \N__44534\,
            I => \N__44453\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__44531\,
            I => \N__44442\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__44528\,
            I => \N__44442\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__44525\,
            I => \N__44442\
        );

    \I__10209\ : Span4Mux_h
    port map (
            O => \N__44520\,
            I => \N__44442\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__44509\,
            I => \N__44442\
        );

    \I__10207\ : Span4Mux_v
    port map (
            O => \N__44506\,
            I => \N__44437\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__44503\,
            I => \N__44437\
        );

    \I__10205\ : Span4Mux_v
    port map (
            O => \N__44500\,
            I => \N__44428\
        );

    \I__10204\ : Span4Mux_v
    port map (
            O => \N__44497\,
            I => \N__44428\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__44492\,
            I => \N__44428\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__44481\,
            I => \N__44428\
        );

    \I__10201\ : CascadeMux
    port map (
            O => \N__44480\,
            I => \N__44414\
        );

    \I__10200\ : CascadeMux
    port map (
            O => \N__44479\,
            I => \N__44409\
        );

    \I__10199\ : InMux
    port map (
            O => \N__44478\,
            I => \N__44401\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44477\,
            I => \N__44401\
        );

    \I__10197\ : InMux
    port map (
            O => \N__44476\,
            I => \N__44401\
        );

    \I__10196\ : Span4Mux_h
    port map (
            O => \N__44471\,
            I => \N__44396\
        );

    \I__10195\ : Span4Mux_v
    port map (
            O => \N__44466\,
            I => \N__44396\
        );

    \I__10194\ : InMux
    port map (
            O => \N__44465\,
            I => \N__44389\
        );

    \I__10193\ : InMux
    port map (
            O => \N__44464\,
            I => \N__44389\
        );

    \I__10192\ : InMux
    port map (
            O => \N__44463\,
            I => \N__44389\
        );

    \I__10191\ : Span4Mux_v
    port map (
            O => \N__44458\,
            I => \N__44386\
        );

    \I__10190\ : InMux
    port map (
            O => \N__44457\,
            I => \N__44381\
        );

    \I__10189\ : InMux
    port map (
            O => \N__44456\,
            I => \N__44381\
        );

    \I__10188\ : LocalMux
    port map (
            O => \N__44453\,
            I => \N__44376\
        );

    \I__10187\ : Span4Mux_v
    port map (
            O => \N__44442\,
            I => \N__44376\
        );

    \I__10186\ : Span4Mux_v
    port map (
            O => \N__44437\,
            I => \N__44371\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__44428\,
            I => \N__44371\
        );

    \I__10184\ : InMux
    port map (
            O => \N__44427\,
            I => \N__44364\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44426\,
            I => \N__44364\
        );

    \I__10182\ : InMux
    port map (
            O => \N__44425\,
            I => \N__44364\
        );

    \I__10181\ : InMux
    port map (
            O => \N__44424\,
            I => \N__44353\
        );

    \I__10180\ : InMux
    port map (
            O => \N__44423\,
            I => \N__44353\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44422\,
            I => \N__44353\
        );

    \I__10178\ : InMux
    port map (
            O => \N__44421\,
            I => \N__44353\
        );

    \I__10177\ : InMux
    port map (
            O => \N__44420\,
            I => \N__44353\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44419\,
            I => \N__44348\
        );

    \I__10175\ : InMux
    port map (
            O => \N__44418\,
            I => \N__44348\
        );

    \I__10174\ : InMux
    port map (
            O => \N__44417\,
            I => \N__44345\
        );

    \I__10173\ : InMux
    port map (
            O => \N__44414\,
            I => \N__44334\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44413\,
            I => \N__44334\
        );

    \I__10171\ : InMux
    port map (
            O => \N__44412\,
            I => \N__44334\
        );

    \I__10170\ : InMux
    port map (
            O => \N__44409\,
            I => \N__44334\
        );

    \I__10169\ : InMux
    port map (
            O => \N__44408\,
            I => \N__44334\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__44401\,
            I => \N__44327\
        );

    \I__10167\ : Span4Mux_h
    port map (
            O => \N__44396\,
            I => \N__44327\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__44389\,
            I => \N__44327\
        );

    \I__10165\ : Odrv4
    port map (
            O => \N__44386\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__44381\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10163\ : Odrv4
    port map (
            O => \N__44376\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10162\ : Odrv4
    port map (
            O => \N__44371\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__44364\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__44353\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__44348\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__44345\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__44334\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10156\ : Odrv4
    port map (
            O => \N__44327\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44306\,
            I => \N__44303\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__44303\,
            I => \N__44300\
        );

    \I__10153\ : Span4Mux_h
    port map (
            O => \N__44300\,
            I => \N__44297\
        );

    \I__10152\ : Odrv4
    port map (
            O => \N__44297\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__10151\ : InMux
    port map (
            O => \N__44294\,
            I => \N__44291\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__44291\,
            I => \N__44288\
        );

    \I__10149\ : Span4Mux_h
    port map (
            O => \N__44288\,
            I => \N__44285\
        );

    \I__10148\ : Odrv4
    port map (
            O => \N__44285\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44282\,
            I => \N__44279\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__44279\,
            I => \N__44276\
        );

    \I__10145\ : Span4Mux_h
    port map (
            O => \N__44276\,
            I => \N__44273\
        );

    \I__10144\ : Odrv4
    port map (
            O => \N__44273\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__10143\ : CascadeMux
    port map (
            O => \N__44270\,
            I => \N__44267\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44267\,
            I => \N__44264\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__44264\,
            I => \N__44261\
        );

    \I__10140\ : Span4Mux_h
    port map (
            O => \N__44261\,
            I => \N__44258\
        );

    \I__10139\ : Odrv4
    port map (
            O => \N__44258\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__10138\ : InMux
    port map (
            O => \N__44255\,
            I => \N__44249\
        );

    \I__10137\ : InMux
    port map (
            O => \N__44254\,
            I => \N__44249\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__44249\,
            I => \N__44246\
        );

    \I__10135\ : Odrv4
    port map (
            O => \N__44246\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__10134\ : CascadeMux
    port map (
            O => \N__44243\,
            I => \N__44239\
        );

    \I__10133\ : CascadeMux
    port map (
            O => \N__44242\,
            I => \N__44236\
        );

    \I__10132\ : InMux
    port map (
            O => \N__44239\,
            I => \N__44233\
        );

    \I__10131\ : InMux
    port map (
            O => \N__44236\,
            I => \N__44230\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__44233\,
            I => \N__44227\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__44230\,
            I => \N__44224\
        );

    \I__10128\ : Span4Mux_v
    port map (
            O => \N__44227\,
            I => \N__44219\
        );

    \I__10127\ : Span4Mux_v
    port map (
            O => \N__44224\,
            I => \N__44219\
        );

    \I__10126\ : Span4Mux_h
    port map (
            O => \N__44219\,
            I => \N__44216\
        );

    \I__10125\ : Odrv4
    port map (
            O => \N__44216\,
            I => \current_shift_inst.un4_control_input_0_31\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44213\,
            I => \N__44210\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__44210\,
            I => \N__44207\
        );

    \I__10122\ : Span4Mux_h
    port map (
            O => \N__44207\,
            I => \N__44204\
        );

    \I__10121\ : Odrv4
    port map (
            O => \N__44204\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44201\,
            I => \N__44198\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__44198\,
            I => \N__44194\
        );

    \I__10118\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44190\
        );

    \I__10117\ : Span4Mux_h
    port map (
            O => \N__44194\,
            I => \N__44187\
        );

    \I__10116\ : InMux
    port map (
            O => \N__44193\,
            I => \N__44184\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__44190\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__10114\ : Odrv4
    port map (
            O => \N__44187\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__44184\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__10112\ : CascadeMux
    port map (
            O => \N__44177\,
            I => \N__44174\
        );

    \I__10111\ : InMux
    port map (
            O => \N__44174\,
            I => \N__44171\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__44171\,
            I => \N__44168\
        );

    \I__10109\ : Odrv12
    port map (
            O => \N__44168\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__10108\ : InMux
    port map (
            O => \N__44165\,
            I => \N__44162\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__44162\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__10106\ : CascadeMux
    port map (
            O => \N__44159\,
            I => \N__44156\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44156\,
            I => \N__44152\
        );

    \I__10104\ : CascadeMux
    port map (
            O => \N__44155\,
            I => \N__44149\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__44152\,
            I => \N__44146\
        );

    \I__10102\ : InMux
    port map (
            O => \N__44149\,
            I => \N__44142\
        );

    \I__10101\ : Span4Mux_h
    port map (
            O => \N__44146\,
            I => \N__44139\
        );

    \I__10100\ : InMux
    port map (
            O => \N__44145\,
            I => \N__44136\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__44142\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10098\ : Odrv4
    port map (
            O => \N__44139\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__44136\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10096\ : InMux
    port map (
            O => \N__44129\,
            I => \N__44126\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__44126\,
            I => \N__44123\
        );

    \I__10094\ : Odrv12
    port map (
            O => \N__44123\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44120\,
            I => \N__44117\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__44117\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__10091\ : CascadeMux
    port map (
            O => \N__44114\,
            I => \N__44111\
        );

    \I__10090\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44108\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44108\,
            I => \N__44105\
        );

    \I__10088\ : Span4Mux_v
    port map (
            O => \N__44105\,
            I => \N__44102\
        );

    \I__10087\ : Odrv4
    port map (
            O => \N__44102\,
            I => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\
        );

    \I__10086\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44095\
        );

    \I__10085\ : CascadeMux
    port map (
            O => \N__44098\,
            I => \N__44089\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__44095\,
            I => \N__44072\
        );

    \I__10083\ : InMux
    port map (
            O => \N__44094\,
            I => \N__44067\
        );

    \I__10082\ : InMux
    port map (
            O => \N__44093\,
            I => \N__44067\
        );

    \I__10081\ : InMux
    port map (
            O => \N__44092\,
            I => \N__44062\
        );

    \I__10080\ : InMux
    port map (
            O => \N__44089\,
            I => \N__44055\
        );

    \I__10079\ : InMux
    port map (
            O => \N__44088\,
            I => \N__44055\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44087\,
            I => \N__44055\
        );

    \I__10077\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44052\
        );

    \I__10076\ : InMux
    port map (
            O => \N__44085\,
            I => \N__44037\
        );

    \I__10075\ : InMux
    port map (
            O => \N__44084\,
            I => \N__44037\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44083\,
            I => \N__44037\
        );

    \I__10073\ : InMux
    port map (
            O => \N__44082\,
            I => \N__44037\
        );

    \I__10072\ : InMux
    port map (
            O => \N__44081\,
            I => \N__44037\
        );

    \I__10071\ : InMux
    port map (
            O => \N__44080\,
            I => \N__44037\
        );

    \I__10070\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44037\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44034\
        );

    \I__10068\ : InMux
    port map (
            O => \N__44077\,
            I => \N__44031\
        );

    \I__10067\ : InMux
    port map (
            O => \N__44076\,
            I => \N__44026\
        );

    \I__10066\ : InMux
    port map (
            O => \N__44075\,
            I => \N__44026\
        );

    \I__10065\ : Span4Mux_v
    port map (
            O => \N__44072\,
            I => \N__44020\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__44067\,
            I => \N__44020\
        );

    \I__10063\ : InMux
    port map (
            O => \N__44066\,
            I => \N__44015\
        );

    \I__10062\ : InMux
    port map (
            O => \N__44065\,
            I => \N__44015\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__44062\,
            I => \N__44007\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__44055\,
            I => \N__44007\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__44052\,
            I => \N__44007\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__44037\,
            I => \N__44004\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__44034\,
            I => \N__44001\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__44031\,
            I => \N__43998\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__44026\,
            I => \N__43993\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44025\,
            I => \N__43990\
        );

    \I__10053\ : Span4Mux_v
    port map (
            O => \N__44020\,
            I => \N__43987\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__44015\,
            I => \N__43984\
        );

    \I__10051\ : InMux
    port map (
            O => \N__44014\,
            I => \N__43981\
        );

    \I__10050\ : Span4Mux_v
    port map (
            O => \N__44007\,
            I => \N__43976\
        );

    \I__10049\ : Span4Mux_v
    port map (
            O => \N__44004\,
            I => \N__43976\
        );

    \I__10048\ : Span4Mux_h
    port map (
            O => \N__44001\,
            I => \N__43973\
        );

    \I__10047\ : Span4Mux_h
    port map (
            O => \N__43998\,
            I => \N__43970\
        );

    \I__10046\ : InMux
    port map (
            O => \N__43997\,
            I => \N__43967\
        );

    \I__10045\ : InMux
    port map (
            O => \N__43996\,
            I => \N__43964\
        );

    \I__10044\ : Span12Mux_h
    port map (
            O => \N__43993\,
            I => \N__43961\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__43990\,
            I => \N__43956\
        );

    \I__10042\ : Span4Mux_h
    port map (
            O => \N__43987\,
            I => \N__43956\
        );

    \I__10041\ : Span4Mux_h
    port map (
            O => \N__43984\,
            I => \N__43947\
        );

    \I__10040\ : LocalMux
    port map (
            O => \N__43981\,
            I => \N__43947\
        );

    \I__10039\ : Span4Mux_h
    port map (
            O => \N__43976\,
            I => \N__43947\
        );

    \I__10038\ : Span4Mux_h
    port map (
            O => \N__43973\,
            I => \N__43947\
        );

    \I__10037\ : Span4Mux_h
    port map (
            O => \N__43970\,
            I => \N__43944\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__43967\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__43964\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10034\ : Odrv12
    port map (
            O => \N__43961\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10033\ : Odrv4
    port map (
            O => \N__43956\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10032\ : Odrv4
    port map (
            O => \N__43947\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10031\ : Odrv4
    port map (
            O => \N__43944\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__10030\ : InMux
    port map (
            O => \N__43931\,
            I => \N__43928\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__43928\,
            I => \N__43924\
        );

    \I__10028\ : InMux
    port map (
            O => \N__43927\,
            I => \N__43920\
        );

    \I__10027\ : Span12Mux_s8_h
    port map (
            O => \N__43924\,
            I => \N__43917\
        );

    \I__10026\ : InMux
    port map (
            O => \N__43923\,
            I => \N__43914\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__43920\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10024\ : Odrv12
    port map (
            O => \N__43917\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__43914\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10022\ : CascadeMux
    port map (
            O => \N__43907\,
            I => \N__43904\
        );

    \I__10021\ : InMux
    port map (
            O => \N__43904\,
            I => \N__43901\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__43901\,
            I => \N__43898\
        );

    \I__10019\ : Odrv12
    port map (
            O => \N__43898\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__10018\ : InMux
    port map (
            O => \N__43895\,
            I => \N__43892\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__43892\,
            I => \N__43889\
        );

    \I__10016\ : Odrv12
    port map (
            O => \N__43889\,
            I => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\
        );

    \I__10015\ : CascadeMux
    port map (
            O => \N__43886\,
            I => \N__43883\
        );

    \I__10014\ : InMux
    port map (
            O => \N__43883\,
            I => \N__43879\
        );

    \I__10013\ : InMux
    port map (
            O => \N__43882\,
            I => \N__43876\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__43879\,
            I => \N__43873\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__43876\,
            I => \N__43869\
        );

    \I__10010\ : Span4Mux_v
    port map (
            O => \N__43873\,
            I => \N__43866\
        );

    \I__10009\ : InMux
    port map (
            O => \N__43872\,
            I => \N__43863\
        );

    \I__10008\ : Odrv12
    port map (
            O => \N__43869\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__10007\ : Odrv4
    port map (
            O => \N__43866\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__43863\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__10005\ : CascadeMux
    port map (
            O => \N__43856\,
            I => \N__43853\
        );

    \I__10004\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43850\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__43850\,
            I => \N__43847\
        );

    \I__10002\ : Span4Mux_h
    port map (
            O => \N__43847\,
            I => \N__43844\
        );

    \I__10001\ : Odrv4
    port map (
            O => \N__43844\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__10000\ : InMux
    port map (
            O => \N__43841\,
            I => \N__43838\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__43838\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__9998\ : CascadeMux
    port map (
            O => \N__43835\,
            I => \N__43832\
        );

    \I__9997\ : InMux
    port map (
            O => \N__43832\,
            I => \N__43829\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__43829\,
            I => \N__43826\
        );

    \I__9995\ : Span4Mux_v
    port map (
            O => \N__43826\,
            I => \N__43823\
        );

    \I__9994\ : Span4Mux_h
    port map (
            O => \N__43823\,
            I => \N__43820\
        );

    \I__9993\ : Odrv4
    port map (
            O => \N__43820\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__9992\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43814\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__43814\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__9990\ : CascadeMux
    port map (
            O => \N__43811\,
            I => \N__43807\
        );

    \I__9989\ : InMux
    port map (
            O => \N__43810\,
            I => \N__43802\
        );

    \I__9988\ : InMux
    port map (
            O => \N__43807\,
            I => \N__43802\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__43802\,
            I => \N__43798\
        );

    \I__9986\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43794\
        );

    \I__9985\ : Span4Mux_h
    port map (
            O => \N__43798\,
            I => \N__43791\
        );

    \I__9984\ : InMux
    port map (
            O => \N__43797\,
            I => \N__43788\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__43794\,
            I => \N__43785\
        );

    \I__9982\ : Odrv4
    port map (
            O => \N__43791\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__43788\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__9980\ : Odrv12
    port map (
            O => \N__43785\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__9979\ : CascadeMux
    port map (
            O => \N__43778\,
            I => \N__43775\
        );

    \I__9978\ : InMux
    port map (
            O => \N__43775\,
            I => \N__43772\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__43772\,
            I => \N__43769\
        );

    \I__9976\ : Span4Mux_v
    port map (
            O => \N__43769\,
            I => \N__43766\
        );

    \I__9975\ : Odrv4
    port map (
            O => \N__43766\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__9974\ : CascadeMux
    port map (
            O => \N__43763\,
            I => \N__43760\
        );

    \I__9973\ : InMux
    port map (
            O => \N__43760\,
            I => \N__43751\
        );

    \I__9972\ : InMux
    port map (
            O => \N__43759\,
            I => \N__43751\
        );

    \I__9971\ : InMux
    port map (
            O => \N__43758\,
            I => \N__43751\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__43751\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__9969\ : InMux
    port map (
            O => \N__43748\,
            I => \N__43736\
        );

    \I__9968\ : InMux
    port map (
            O => \N__43747\,
            I => \N__43736\
        );

    \I__9967\ : InMux
    port map (
            O => \N__43746\,
            I => \N__43736\
        );

    \I__9966\ : InMux
    port map (
            O => \N__43745\,
            I => \N__43736\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__43736\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__9964\ : CascadeMux
    port map (
            O => \N__43733\,
            I => \N__43730\
        );

    \I__9963\ : InMux
    port map (
            O => \N__43730\,
            I => \N__43727\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__43727\,
            I => \N__43724\
        );

    \I__9961\ : Span4Mux_h
    port map (
            O => \N__43724\,
            I => \N__43721\
        );

    \I__9960\ : Odrv4
    port map (
            O => \N__43721\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__9959\ : InMux
    port map (
            O => \N__43718\,
            I => \N__43715\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__43715\,
            I => \N__43712\
        );

    \I__9957\ : Odrv4
    port map (
            O => \N__43712\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__9956\ : InMux
    port map (
            O => \N__43709\,
            I => \N__43705\
        );

    \I__9955\ : CascadeMux
    port map (
            O => \N__43708\,
            I => \N__43702\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__43705\,
            I => \N__43698\
        );

    \I__9953\ : InMux
    port map (
            O => \N__43702\,
            I => \N__43693\
        );

    \I__9952\ : InMux
    port map (
            O => \N__43701\,
            I => \N__43693\
        );

    \I__9951\ : Span4Mux_v
    port map (
            O => \N__43698\,
            I => \N__43690\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__43693\,
            I => \N__43687\
        );

    \I__9949\ : Odrv4
    port map (
            O => \N__43690\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9948\ : Odrv4
    port map (
            O => \N__43687\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9947\ : CascadeMux
    port map (
            O => \N__43682\,
            I => \N__43679\
        );

    \I__9946\ : InMux
    port map (
            O => \N__43679\,
            I => \N__43676\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__43676\,
            I => \N__43673\
        );

    \I__9944\ : Span4Mux_v
    port map (
            O => \N__43673\,
            I => \N__43670\
        );

    \I__9943\ : Odrv4
    port map (
            O => \N__43670\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__9942\ : CascadeMux
    port map (
            O => \N__43667\,
            I => \N__43664\
        );

    \I__9941\ : InMux
    port map (
            O => \N__43664\,
            I => \N__43660\
        );

    \I__9940\ : CascadeMux
    port map (
            O => \N__43663\,
            I => \N__43657\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__43660\,
            I => \N__43654\
        );

    \I__9938\ : InMux
    port map (
            O => \N__43657\,
            I => \N__43651\
        );

    \I__9937\ : Span4Mux_v
    port map (
            O => \N__43654\,
            I => \N__43647\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__43651\,
            I => \N__43644\
        );

    \I__9935\ : InMux
    port map (
            O => \N__43650\,
            I => \N__43641\
        );

    \I__9934\ : Span4Mux_h
    port map (
            O => \N__43647\,
            I => \N__43638\
        );

    \I__9933\ : Span4Mux_h
    port map (
            O => \N__43644\,
            I => \N__43635\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__43641\,
            I => \N__43632\
        );

    \I__9931\ : Odrv4
    port map (
            O => \N__43638\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9930\ : Odrv4
    port map (
            O => \N__43635\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9929\ : Odrv4
    port map (
            O => \N__43632\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9928\ : InMux
    port map (
            O => \N__43625\,
            I => \N__43622\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__43622\,
            I => \N__43619\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__43619\,
            I => \N__43616\
        );

    \I__9925\ : Odrv4
    port map (
            O => \N__43616\,
            I => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\
        );

    \I__9924\ : InMux
    port map (
            O => \N__43613\,
            I => \N__43608\
        );

    \I__9923\ : InMux
    port map (
            O => \N__43612\,
            I => \N__43605\
        );

    \I__9922\ : InMux
    port map (
            O => \N__43611\,
            I => \N__43602\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__43608\,
            I => \N__43599\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__43605\,
            I => \N__43596\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__43602\,
            I => \N__43593\
        );

    \I__9918\ : Odrv12
    port map (
            O => \N__43599\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__43596\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9916\ : Odrv4
    port map (
            O => \N__43593\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9915\ : CascadeMux
    port map (
            O => \N__43586\,
            I => \N__43583\
        );

    \I__9914\ : InMux
    port map (
            O => \N__43583\,
            I => \N__43580\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__43580\,
            I => \N__43577\
        );

    \I__9912\ : Span4Mux_v
    port map (
            O => \N__43577\,
            I => \N__43574\
        );

    \I__9911\ : Span4Mux_h
    port map (
            O => \N__43574\,
            I => \N__43571\
        );

    \I__9910\ : Odrv4
    port map (
            O => \N__43571\,
            I => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\
        );

    \I__9909\ : CascadeMux
    port map (
            O => \N__43568\,
            I => \N__43565\
        );

    \I__9908\ : InMux
    port map (
            O => \N__43565\,
            I => \N__43562\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__43562\,
            I => \N__43559\
        );

    \I__9906\ : Span4Mux_v
    port map (
            O => \N__43559\,
            I => \N__43556\
        );

    \I__9905\ : Odrv4
    port map (
            O => \N__43556\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__9904\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43549\
        );

    \I__9903\ : InMux
    port map (
            O => \N__43552\,
            I => \N__43546\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__43549\,
            I => \N__43542\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__43546\,
            I => \N__43539\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43545\,
            I => \N__43536\
        );

    \I__9899\ : Span4Mux_v
    port map (
            O => \N__43542\,
            I => \N__43533\
        );

    \I__9898\ : Odrv12
    port map (
            O => \N__43539\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__43536\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9896\ : Odrv4
    port map (
            O => \N__43533\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9895\ : CascadeMux
    port map (
            O => \N__43526\,
            I => \N__43523\
        );

    \I__9894\ : InMux
    port map (
            O => \N__43523\,
            I => \N__43520\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__43520\,
            I => \N__43517\
        );

    \I__9892\ : Span4Mux_h
    port map (
            O => \N__43517\,
            I => \N__43514\
        );

    \I__9891\ : Span4Mux_v
    port map (
            O => \N__43514\,
            I => \N__43511\
        );

    \I__9890\ : Odrv4
    port map (
            O => \N__43511\,
            I => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\
        );

    \I__9889\ : CascadeMux
    port map (
            O => \N__43508\,
            I => \N__43505\
        );

    \I__9888\ : InMux
    port map (
            O => \N__43505\,
            I => \N__43501\
        );

    \I__9887\ : InMux
    port map (
            O => \N__43504\,
            I => \N__43498\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__43501\,
            I => \N__43494\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__43498\,
            I => \N__43491\
        );

    \I__9884\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43488\
        );

    \I__9883\ : Span4Mux_v
    port map (
            O => \N__43494\,
            I => \N__43483\
        );

    \I__9882\ : Span4Mux_v
    port map (
            O => \N__43491\,
            I => \N__43483\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__43488\,
            I => \N__43480\
        );

    \I__9880\ : Odrv4
    port map (
            O => \N__43483\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9879\ : Odrv4
    port map (
            O => \N__43480\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9878\ : CascadeMux
    port map (
            O => \N__43475\,
            I => \N__43472\
        );

    \I__9877\ : InMux
    port map (
            O => \N__43472\,
            I => \N__43469\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__43469\,
            I => \N__43466\
        );

    \I__9875\ : Span4Mux_h
    port map (
            O => \N__43466\,
            I => \N__43463\
        );

    \I__9874\ : Odrv4
    port map (
            O => \N__43463\,
            I => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43460\,
            I => \N__43457\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__43457\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__9871\ : InMux
    port map (
            O => \N__43454\,
            I => \N__43451\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__43451\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__9869\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43444\
        );

    \I__9868\ : InMux
    port map (
            O => \N__43447\,
            I => \N__43441\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__43444\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__43441\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9865\ : InMux
    port map (
            O => \N__43436\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__9864\ : InMux
    port map (
            O => \N__43433\,
            I => \N__43429\
        );

    \I__9863\ : InMux
    port map (
            O => \N__43432\,
            I => \N__43426\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__43429\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__43426\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9860\ : InMux
    port map (
            O => \N__43421\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__9859\ : InMux
    port map (
            O => \N__43418\,
            I => \N__43414\
        );

    \I__9858\ : InMux
    port map (
            O => \N__43417\,
            I => \N__43411\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__43414\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__43411\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9855\ : InMux
    port map (
            O => \N__43406\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43403\,
            I => \N__43399\
        );

    \I__9853\ : InMux
    port map (
            O => \N__43402\,
            I => \N__43396\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__43399\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__43396\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43391\,
            I => \bfn_18_13_0_\
        );

    \I__9849\ : InMux
    port map (
            O => \N__43388\,
            I => \N__43384\
        );

    \I__9848\ : InMux
    port map (
            O => \N__43387\,
            I => \N__43381\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__43384\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__43381\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9845\ : InMux
    port map (
            O => \N__43376\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__9844\ : CEMux
    port map (
            O => \N__43373\,
            I => \N__43364\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43372\,
            I => \N__43355\
        );

    \I__9842\ : InMux
    port map (
            O => \N__43371\,
            I => \N__43355\
        );

    \I__9841\ : InMux
    port map (
            O => \N__43370\,
            I => \N__43355\
        );

    \I__9840\ : InMux
    port map (
            O => \N__43369\,
            I => \N__43355\
        );

    \I__9839\ : CEMux
    port map (
            O => \N__43368\,
            I => \N__43352\
        );

    \I__9838\ : CEMux
    port map (
            O => \N__43367\,
            I => \N__43348\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__43364\,
            I => \N__43345\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__43355\,
            I => \N__43340\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__43352\,
            I => \N__43340\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43351\,
            I => \N__43323\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__43348\,
            I => \N__43318\
        );

    \I__9832\ : Span4Mux_h
    port map (
            O => \N__43345\,
            I => \N__43318\
        );

    \I__9831\ : Span4Mux_v
    port map (
            O => \N__43340\,
            I => \N__43315\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43339\,
            I => \N__43308\
        );

    \I__9829\ : InMux
    port map (
            O => \N__43338\,
            I => \N__43308\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43337\,
            I => \N__43308\
        );

    \I__9827\ : InMux
    port map (
            O => \N__43336\,
            I => \N__43299\
        );

    \I__9826\ : InMux
    port map (
            O => \N__43335\,
            I => \N__43299\
        );

    \I__9825\ : InMux
    port map (
            O => \N__43334\,
            I => \N__43299\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43333\,
            I => \N__43299\
        );

    \I__9823\ : InMux
    port map (
            O => \N__43332\,
            I => \N__43296\
        );

    \I__9822\ : InMux
    port map (
            O => \N__43331\,
            I => \N__43291\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43330\,
            I => \N__43291\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43329\,
            I => \N__43282\
        );

    \I__9819\ : InMux
    port map (
            O => \N__43328\,
            I => \N__43282\
        );

    \I__9818\ : InMux
    port map (
            O => \N__43327\,
            I => \N__43282\
        );

    \I__9817\ : InMux
    port map (
            O => \N__43326\,
            I => \N__43282\
        );

    \I__9816\ : LocalMux
    port map (
            O => \N__43323\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__9815\ : Odrv4
    port map (
            O => \N__43318\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__9814\ : Odrv4
    port map (
            O => \N__43315\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__43308\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__43299\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__43296\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43291\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__43282\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__9808\ : InMux
    port map (
            O => \N__43265\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__9807\ : InMux
    port map (
            O => \N__43262\,
            I => \N__43258\
        );

    \I__9806\ : InMux
    port map (
            O => \N__43261\,
            I => \N__43255\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__43258\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__43255\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9803\ : InMux
    port map (
            O => \N__43250\,
            I => \N__43245\
        );

    \I__9802\ : InMux
    port map (
            O => \N__43249\,
            I => \N__43242\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43248\,
            I => \N__43239\
        );

    \I__9800\ : LocalMux
    port map (
            O => \N__43245\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__43242\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__43239\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9797\ : CascadeMux
    port map (
            O => \N__43232\,
            I => \N__43229\
        );

    \I__9796\ : InMux
    port map (
            O => \N__43229\,
            I => \N__43226\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__43226\,
            I => \N__43223\
        );

    \I__9794\ : Span4Mux_h
    port map (
            O => \N__43223\,
            I => \N__43220\
        );

    \I__9793\ : Span4Mux_v
    port map (
            O => \N__43220\,
            I => \N__43217\
        );

    \I__9792\ : Odrv4
    port map (
            O => \N__43217\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__9791\ : CascadeMux
    port map (
            O => \N__43214\,
            I => \N__43211\
        );

    \I__9790\ : InMux
    port map (
            O => \N__43211\,
            I => \N__43208\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__43208\,
            I => \N__43205\
        );

    \I__9788\ : Span4Mux_h
    port map (
            O => \N__43205\,
            I => \N__43202\
        );

    \I__9787\ : Odrv4
    port map (
            O => \N__43202\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__9786\ : CascadeMux
    port map (
            O => \N__43199\,
            I => \N__43196\
        );

    \I__9785\ : InMux
    port map (
            O => \N__43196\,
            I => \N__43193\
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__43193\,
            I => \N__43190\
        );

    \I__9783\ : Span4Mux_v
    port map (
            O => \N__43190\,
            I => \N__43187\
        );

    \I__9782\ : Span4Mux_h
    port map (
            O => \N__43187\,
            I => \N__43184\
        );

    \I__9781\ : Odrv4
    port map (
            O => \N__43184\,
            I => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\
        );

    \I__9780\ : InMux
    port map (
            O => \N__43181\,
            I => \N__43177\
        );

    \I__9779\ : InMux
    port map (
            O => \N__43180\,
            I => \N__43174\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__43177\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__43174\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__9776\ : InMux
    port map (
            O => \N__43169\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__9775\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43162\
        );

    \I__9774\ : InMux
    port map (
            O => \N__43165\,
            I => \N__43159\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__43162\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__43159\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9771\ : InMux
    port map (
            O => \N__43154\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43151\,
            I => \N__43147\
        );

    \I__9769\ : InMux
    port map (
            O => \N__43150\,
            I => \N__43144\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__43147\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__43144\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43139\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__9765\ : InMux
    port map (
            O => \N__43136\,
            I => \N__43132\
        );

    \I__9764\ : InMux
    port map (
            O => \N__43135\,
            I => \N__43129\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__43132\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__43129\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__9761\ : InMux
    port map (
            O => \N__43124\,
            I => \bfn_18_12_0_\
        );

    \I__9760\ : InMux
    port map (
            O => \N__43121\,
            I => \N__43117\
        );

    \I__9759\ : InMux
    port map (
            O => \N__43120\,
            I => \N__43114\
        );

    \I__9758\ : LocalMux
    port map (
            O => \N__43117\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__43114\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__9756\ : InMux
    port map (
            O => \N__43109\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__9755\ : InMux
    port map (
            O => \N__43106\,
            I => \N__43102\
        );

    \I__9754\ : InMux
    port map (
            O => \N__43105\,
            I => \N__43099\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__43102\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__43099\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__9751\ : InMux
    port map (
            O => \N__43094\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__9750\ : InMux
    port map (
            O => \N__43091\,
            I => \N__43087\
        );

    \I__9749\ : InMux
    port map (
            O => \N__43090\,
            I => \N__43084\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__43087\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__43084\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__9746\ : InMux
    port map (
            O => \N__43079\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__9745\ : InMux
    port map (
            O => \N__43076\,
            I => \N__43072\
        );

    \I__9744\ : InMux
    port map (
            O => \N__43075\,
            I => \N__43069\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__43072\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__43069\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__9741\ : InMux
    port map (
            O => \N__43064\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__9740\ : InMux
    port map (
            O => \N__43061\,
            I => \N__43058\
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__43058\,
            I => \N__43055\
        );

    \I__9738\ : Span4Mux_v
    port map (
            O => \N__43055\,
            I => \N__43051\
        );

    \I__9737\ : InMux
    port map (
            O => \N__43054\,
            I => \N__43048\
        );

    \I__9736\ : Odrv4
    port map (
            O => \N__43051\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__43048\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__9734\ : InMux
    port map (
            O => \N__43043\,
            I => \N__43040\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__43040\,
            I => \N__43037\
        );

    \I__9732\ : Span12Mux_h
    port map (
            O => \N__43037\,
            I => \N__43034\
        );

    \I__9731\ : Odrv12
    port map (
            O => \N__43034\,
            I => \phase_controller_inst1.stoper_tr.running_1_sqmuxa\
        );

    \I__9730\ : InMux
    port map (
            O => \N__43031\,
            I => \N__43025\
        );

    \I__9729\ : InMux
    port map (
            O => \N__43030\,
            I => \N__43025\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__43025\,
            I => \N__43017\
        );

    \I__9727\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43013\
        );

    \I__9726\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43010\
        );

    \I__9725\ : InMux
    port map (
            O => \N__43022\,
            I => \N__43005\
        );

    \I__9724\ : InMux
    port map (
            O => \N__43021\,
            I => \N__43005\
        );

    \I__9723\ : InMux
    port map (
            O => \N__43020\,
            I => \N__43002\
        );

    \I__9722\ : Span4Mux_h
    port map (
            O => \N__43017\,
            I => \N__42999\
        );

    \I__9721\ : InMux
    port map (
            O => \N__43016\,
            I => \N__42996\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__43013\,
            I => \N__42989\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__43010\,
            I => \N__42989\
        );

    \I__9718\ : LocalMux
    port map (
            O => \N__43005\,
            I => \N__42989\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__43002\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9716\ : Odrv4
    port map (
            O => \N__42999\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__42996\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9714\ : Odrv12
    port map (
            O => \N__42989\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9713\ : CascadeMux
    port map (
            O => \N__42980\,
            I => \N__42976\
        );

    \I__9712\ : InMux
    port map (
            O => \N__42979\,
            I => \N__42972\
        );

    \I__9711\ : InMux
    port map (
            O => \N__42976\,
            I => \N__42968\
        );

    \I__9710\ : CascadeMux
    port map (
            O => \N__42975\,
            I => \N__42965\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__42972\,
            I => \N__42962\
        );

    \I__9708\ : InMux
    port map (
            O => \N__42971\,
            I => \N__42959\
        );

    \I__9707\ : LocalMux
    port map (
            O => \N__42968\,
            I => \N__42955\
        );

    \I__9706\ : InMux
    port map (
            O => \N__42965\,
            I => \N__42952\
        );

    \I__9705\ : Span4Mux_v
    port map (
            O => \N__42962\,
            I => \N__42949\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__42959\,
            I => \N__42946\
        );

    \I__9703\ : InMux
    port map (
            O => \N__42958\,
            I => \N__42941\
        );

    \I__9702\ : Span4Mux_h
    port map (
            O => \N__42955\,
            I => \N__42938\
        );

    \I__9701\ : LocalMux
    port map (
            O => \N__42952\,
            I => \N__42931\
        );

    \I__9700\ : Span4Mux_h
    port map (
            O => \N__42949\,
            I => \N__42931\
        );

    \I__9699\ : Span4Mux_v
    port map (
            O => \N__42946\,
            I => \N__42931\
        );

    \I__9698\ : InMux
    port map (
            O => \N__42945\,
            I => \N__42926\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42944\,
            I => \N__42926\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__42941\,
            I => \N__42923\
        );

    \I__9695\ : Odrv4
    port map (
            O => \N__42938\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__9694\ : Odrv4
    port map (
            O => \N__42931\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__42926\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__9692\ : Odrv12
    port map (
            O => \N__42923\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__9691\ : CascadeMux
    port map (
            O => \N__42914\,
            I => \phase_controller_inst1.stoper_tr.running_1_sqmuxa_cascade_\
        );

    \I__9690\ : InMux
    port map (
            O => \N__42911\,
            I => \N__42908\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__42908\,
            I => \N__42904\
        );

    \I__9688\ : InMux
    port map (
            O => \N__42907\,
            I => \N__42901\
        );

    \I__9687\ : Span4Mux_h
    port map (
            O => \N__42904\,
            I => \N__42897\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__42901\,
            I => \N__42894\
        );

    \I__9685\ : InMux
    port map (
            O => \N__42900\,
            I => \N__42891\
        );

    \I__9684\ : Span4Mux_h
    port map (
            O => \N__42897\,
            I => \N__42888\
        );

    \I__9683\ : Span4Mux_h
    port map (
            O => \N__42894\,
            I => \N__42885\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__42891\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__9681\ : Odrv4
    port map (
            O => \N__42888\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__9680\ : Odrv4
    port map (
            O => \N__42885\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__9679\ : InMux
    port map (
            O => \N__42878\,
            I => \N__42875\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__42875\,
            I => \N__42872\
        );

    \I__9677\ : Span4Mux_h
    port map (
            O => \N__42872\,
            I => \N__42869\
        );

    \I__9676\ : Odrv4
    port map (
            O => \N__42869\,
            I => \phase_controller_inst1.stoper_tr.un1_start_latched2_0\
        );

    \I__9675\ : InMux
    port map (
            O => \N__42866\,
            I => \N__42861\
        );

    \I__9674\ : InMux
    port map (
            O => \N__42865\,
            I => \N__42858\
        );

    \I__9673\ : InMux
    port map (
            O => \N__42864\,
            I => \N__42855\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__42861\,
            I => \N__42852\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__42858\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__42855\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__9669\ : Odrv4
    port map (
            O => \N__42852\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42845\,
            I => \N__42841\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42844\,
            I => \N__42836\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__42841\,
            I => \N__42833\
        );

    \I__9665\ : InMux
    port map (
            O => \N__42840\,
            I => \N__42830\
        );

    \I__9664\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42827\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__42836\,
            I => \N__42824\
        );

    \I__9662\ : Span4Mux_v
    port map (
            O => \N__42833\,
            I => \N__42821\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__42830\,
            I => \N__42816\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__42827\,
            I => \N__42816\
        );

    \I__9659\ : Span4Mux_h
    port map (
            O => \N__42824\,
            I => \N__42813\
        );

    \I__9658\ : Odrv4
    port map (
            O => \N__42821\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9657\ : Odrv12
    port map (
            O => \N__42816\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9656\ : Odrv4
    port map (
            O => \N__42813\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__9655\ : InMux
    port map (
            O => \N__42806\,
            I => \N__42803\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__42803\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__9653\ : CascadeMux
    port map (
            O => \N__42800\,
            I => \N__42797\
        );

    \I__9652\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42792\
        );

    \I__9651\ : InMux
    port map (
            O => \N__42796\,
            I => \N__42789\
        );

    \I__9650\ : CascadeMux
    port map (
            O => \N__42795\,
            I => \N__42786\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__42792\,
            I => \N__42783\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__42789\,
            I => \N__42780\
        );

    \I__9647\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42777\
        );

    \I__9646\ : Span4Mux_h
    port map (
            O => \N__42783\,
            I => \N__42774\
        );

    \I__9645\ : Span4Mux_v
    port map (
            O => \N__42780\,
            I => \N__42771\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__42777\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__9643\ : Odrv4
    port map (
            O => \N__42774\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__9642\ : Odrv4
    port map (
            O => \N__42771\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__9641\ : InMux
    port map (
            O => \N__42764\,
            I => \N__42760\
        );

    \I__9640\ : InMux
    port map (
            O => \N__42763\,
            I => \N__42757\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__42760\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__42757\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__9637\ : InMux
    port map (
            O => \N__42752\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__9636\ : InMux
    port map (
            O => \N__42749\,
            I => \N__42746\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__42746\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8IZ0Z2\
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__42743\,
            I => \N__42740\
        );

    \I__9633\ : InMux
    port map (
            O => \N__42740\,
            I => \N__42736\
        );

    \I__9632\ : InMux
    port map (
            O => \N__42739\,
            I => \N__42733\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__42736\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__42733\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__9629\ : InMux
    port map (
            O => \N__42728\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__9628\ : InMux
    port map (
            O => \N__42725\,
            I => \N__42721\
        );

    \I__9627\ : InMux
    port map (
            O => \N__42724\,
            I => \N__42718\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__42721\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__42718\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42713\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__9623\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42706\
        );

    \I__9622\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42703\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__42706\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__42703\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__9619\ : InMux
    port map (
            O => \N__42698\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__9618\ : InMux
    port map (
            O => \N__42695\,
            I => \N__42692\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__42692\,
            I => \N__42687\
        );

    \I__9616\ : InMux
    port map (
            O => \N__42691\,
            I => \N__42684\
        );

    \I__9615\ : InMux
    port map (
            O => \N__42690\,
            I => \N__42681\
        );

    \I__9614\ : Span4Mux_h
    port map (
            O => \N__42687\,
            I => \N__42678\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__42684\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__42681\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6\
        );

    \I__9611\ : Odrv4
    port map (
            O => \N__42678\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6\
        );

    \I__9610\ : CascadeMux
    port map (
            O => \N__42671\,
            I => \N__42668\
        );

    \I__9609\ : InMux
    port map (
            O => \N__42668\,
            I => \N__42665\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__42665\,
            I => \phase_controller_inst1.stoper_tr.un6_running_6\
        );

    \I__9607\ : InMux
    port map (
            O => \N__42662\,
            I => \N__42658\
        );

    \I__9606\ : InMux
    port map (
            O => \N__42661\,
            I => \N__42655\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__42658\,
            I => \N__42652\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__42655\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\
        );

    \I__9603\ : Odrv12
    port map (
            O => \N__42652\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\
        );

    \I__9602\ : InMux
    port map (
            O => \N__42647\,
            I => \N__42644\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__42644\,
            I => \phase_controller_inst1.stoper_tr.un6_running_2\
        );

    \I__9600\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42638\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__42638\,
            I => \phase_controller_inst1.stoper_tr.un6_running_4\
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__42635\,
            I => \N__42632\
        );

    \I__9597\ : InMux
    port map (
            O => \N__42632\,
            I => \N__42629\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__42629\,
            I => \phase_controller_inst1.stoper_tr.un6_running_5\
        );

    \I__9595\ : CascadeMux
    port map (
            O => \N__42626\,
            I => \N__42622\
        );

    \I__9594\ : InMux
    port map (
            O => \N__42625\,
            I => \N__42618\
        );

    \I__9593\ : InMux
    port map (
            O => \N__42622\,
            I => \N__42615\
        );

    \I__9592\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42611\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__42618\,
            I => \N__42608\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__42615\,
            I => \N__42605\
        );

    \I__9589\ : InMux
    port map (
            O => \N__42614\,
            I => \N__42602\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__42611\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__9587\ : Odrv12
    port map (
            O => \N__42608\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__9586\ : Odrv4
    port map (
            O => \N__42605\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__42602\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__9584\ : InMux
    port map (
            O => \N__42593\,
            I => \N__42590\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__42590\,
            I => \phase_controller_inst1.stoper_tr.un6_running_7\
        );

    \I__9582\ : CascadeMux
    port map (
            O => \N__42587\,
            I => \N__42583\
        );

    \I__9581\ : CascadeMux
    port map (
            O => \N__42586\,
            I => \N__42580\
        );

    \I__9580\ : InMux
    port map (
            O => \N__42583\,
            I => \N__42577\
        );

    \I__9579\ : InMux
    port map (
            O => \N__42580\,
            I => \N__42574\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__42577\,
            I => \N__42571\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__42574\,
            I => \N__42568\
        );

    \I__9576\ : Span4Mux_h
    port map (
            O => \N__42571\,
            I => \N__42564\
        );

    \I__9575\ : Span4Mux_h
    port map (
            O => \N__42568\,
            I => \N__42561\
        );

    \I__9574\ : InMux
    port map (
            O => \N__42567\,
            I => \N__42558\
        );

    \I__9573\ : Odrv4
    port map (
            O => \N__42564\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__9572\ : Odrv4
    port map (
            O => \N__42561\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__42558\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__9570\ : CascadeMux
    port map (
            O => \N__42551\,
            I => \N__42548\
        );

    \I__9569\ : InMux
    port map (
            O => \N__42548\,
            I => \N__42545\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__42545\,
            I => \N__42542\
        );

    \I__9567\ : Span4Mux_h
    port map (
            O => \N__42542\,
            I => \N__42539\
        );

    \I__9566\ : Odrv4
    port map (
            O => \N__42539\,
            I => \phase_controller_inst2.stoper_tr.un6_running_4\
        );

    \I__9565\ : InMux
    port map (
            O => \N__42536\,
            I => \N__42499\
        );

    \I__9564\ : InMux
    port map (
            O => \N__42535\,
            I => \N__42499\
        );

    \I__9563\ : InMux
    port map (
            O => \N__42534\,
            I => \N__42499\
        );

    \I__9562\ : InMux
    port map (
            O => \N__42533\,
            I => \N__42499\
        );

    \I__9561\ : InMux
    port map (
            O => \N__42532\,
            I => \N__42499\
        );

    \I__9560\ : InMux
    port map (
            O => \N__42531\,
            I => \N__42494\
        );

    \I__9559\ : InMux
    port map (
            O => \N__42530\,
            I => \N__42494\
        );

    \I__9558\ : InMux
    port map (
            O => \N__42529\,
            I => \N__42479\
        );

    \I__9557\ : InMux
    port map (
            O => \N__42528\,
            I => \N__42479\
        );

    \I__9556\ : InMux
    port map (
            O => \N__42527\,
            I => \N__42479\
        );

    \I__9555\ : InMux
    port map (
            O => \N__42526\,
            I => \N__42479\
        );

    \I__9554\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42479\
        );

    \I__9553\ : InMux
    port map (
            O => \N__42524\,
            I => \N__42479\
        );

    \I__9552\ : InMux
    port map (
            O => \N__42523\,
            I => \N__42479\
        );

    \I__9551\ : InMux
    port map (
            O => \N__42522\,
            I => \N__42468\
        );

    \I__9550\ : InMux
    port map (
            O => \N__42521\,
            I => \N__42468\
        );

    \I__9549\ : InMux
    port map (
            O => \N__42520\,
            I => \N__42468\
        );

    \I__9548\ : InMux
    port map (
            O => \N__42519\,
            I => \N__42468\
        );

    \I__9547\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42468\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42454\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42516\,
            I => \N__42454\
        );

    \I__9544\ : InMux
    port map (
            O => \N__42515\,
            I => \N__42454\
        );

    \I__9543\ : InMux
    port map (
            O => \N__42514\,
            I => \N__42454\
        );

    \I__9542\ : InMux
    port map (
            O => \N__42513\,
            I => \N__42454\
        );

    \I__9541\ : InMux
    port map (
            O => \N__42512\,
            I => \N__42454\
        );

    \I__9540\ : InMux
    port map (
            O => \N__42511\,
            I => \N__42445\
        );

    \I__9539\ : InMux
    port map (
            O => \N__42510\,
            I => \N__42445\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__42499\,
            I => \N__42442\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__42494\,
            I => \N__42439\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__42479\,
            I => \N__42434\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__42468\,
            I => \N__42434\
        );

    \I__9534\ : InMux
    port map (
            O => \N__42467\,
            I => \N__42428\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__42454\,
            I => \N__42425\
        );

    \I__9532\ : InMux
    port map (
            O => \N__42453\,
            I => \N__42422\
        );

    \I__9531\ : InMux
    port map (
            O => \N__42452\,
            I => \N__42419\
        );

    \I__9530\ : InMux
    port map (
            O => \N__42451\,
            I => \N__42414\
        );

    \I__9529\ : InMux
    port map (
            O => \N__42450\,
            I => \N__42414\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__42445\,
            I => \N__42409\
        );

    \I__9527\ : Span4Mux_h
    port map (
            O => \N__42442\,
            I => \N__42409\
        );

    \I__9526\ : Span4Mux_h
    port map (
            O => \N__42439\,
            I => \N__42404\
        );

    \I__9525\ : Span4Mux_v
    port map (
            O => \N__42434\,
            I => \N__42404\
        );

    \I__9524\ : InMux
    port map (
            O => \N__42433\,
            I => \N__42397\
        );

    \I__9523\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42397\
        );

    \I__9522\ : InMux
    port map (
            O => \N__42431\,
            I => \N__42397\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__42428\,
            I => \N__42388\
        );

    \I__9520\ : Span4Mux_v
    port map (
            O => \N__42425\,
            I => \N__42388\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__42422\,
            I => \N__42388\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__42419\,
            I => \N__42388\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__42414\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9516\ : Odrv4
    port map (
            O => \N__42409\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9515\ : Odrv4
    port map (
            O => \N__42404\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__42397\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9513\ : Odrv4
    port map (
            O => \N__42388\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9512\ : InMux
    port map (
            O => \N__42377\,
            I => \N__42374\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__42374\,
            I => \N__42370\
        );

    \I__9510\ : InMux
    port map (
            O => \N__42373\,
            I => \N__42367\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__42370\,
            I => \N__42361\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__42367\,
            I => \N__42361\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42366\,
            I => \N__42357\
        );

    \I__9506\ : Span4Mux_h
    port map (
            O => \N__42361\,
            I => \N__42354\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42360\,
            I => \N__42351\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__42357\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__9503\ : Odrv4
    port map (
            O => \N__42354\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__42351\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__9501\ : InMux
    port map (
            O => \N__42344\,
            I => \N__42341\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__42341\,
            I => \N__42338\
        );

    \I__9499\ : Span4Mux_h
    port map (
            O => \N__42338\,
            I => \N__42335\
        );

    \I__9498\ : Odrv4
    port map (
            O => \N__42335\,
            I => \phase_controller_inst2.stoper_tr.un6_running_5\
        );

    \I__9497\ : CascadeMux
    port map (
            O => \N__42332\,
            I => \N__42328\
        );

    \I__9496\ : InMux
    port map (
            O => \N__42331\,
            I => \N__42325\
        );

    \I__9495\ : InMux
    port map (
            O => \N__42328\,
            I => \N__42322\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42325\,
            I => \N__42319\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__42322\,
            I => \N__42316\
        );

    \I__9492\ : Span4Mux_h
    port map (
            O => \N__42319\,
            I => \N__42313\
        );

    \I__9491\ : Odrv12
    port map (
            O => \N__42316\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\
        );

    \I__9490\ : Odrv4
    port map (
            O => \N__42313\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\
        );

    \I__9489\ : CascadeMux
    port map (
            O => \N__42308\,
            I => \N__42300\
        );

    \I__9488\ : CascadeMux
    port map (
            O => \N__42307\,
            I => \N__42297\
        );

    \I__9487\ : InMux
    port map (
            O => \N__42306\,
            I => \N__42282\
        );

    \I__9486\ : InMux
    port map (
            O => \N__42305\,
            I => \N__42282\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42304\,
            I => \N__42282\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42303\,
            I => \N__42279\
        );

    \I__9483\ : InMux
    port map (
            O => \N__42300\,
            I => \N__42268\
        );

    \I__9482\ : InMux
    port map (
            O => \N__42297\,
            I => \N__42268\
        );

    \I__9481\ : InMux
    port map (
            O => \N__42296\,
            I => \N__42268\
        );

    \I__9480\ : InMux
    port map (
            O => \N__42295\,
            I => \N__42268\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42268\
        );

    \I__9478\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42261\
        );

    \I__9477\ : InMux
    port map (
            O => \N__42292\,
            I => \N__42261\
        );

    \I__9476\ : InMux
    port map (
            O => \N__42291\,
            I => \N__42261\
        );

    \I__9475\ : InMux
    port map (
            O => \N__42290\,
            I => \N__42256\
        );

    \I__9474\ : InMux
    port map (
            O => \N__42289\,
            I => \N__42256\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__42282\,
            I => \N__42253\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__42279\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42268\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__42261\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__42256\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6\
        );

    \I__9468\ : Odrv4
    port map (
            O => \N__42253\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6\
        );

    \I__9467\ : CascadeMux
    port map (
            O => \N__42242\,
            I => \N__42236\
        );

    \I__9466\ : CascadeMux
    port map (
            O => \N__42241\,
            I => \N__42233\
        );

    \I__9465\ : CascadeMux
    port map (
            O => \N__42240\,
            I => \N__42228\
        );

    \I__9464\ : CascadeMux
    port map (
            O => \N__42239\,
            I => \N__42225\
        );

    \I__9463\ : InMux
    port map (
            O => \N__42236\,
            I => \N__42217\
        );

    \I__9462\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42212\
        );

    \I__9461\ : InMux
    port map (
            O => \N__42232\,
            I => \N__42212\
        );

    \I__9460\ : InMux
    port map (
            O => \N__42231\,
            I => \N__42209\
        );

    \I__9459\ : InMux
    port map (
            O => \N__42228\,
            I => \N__42206\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42225\,
            I => \N__42203\
        );

    \I__9457\ : InMux
    port map (
            O => \N__42224\,
            I => \N__42200\
        );

    \I__9456\ : InMux
    port map (
            O => \N__42223\,
            I => \N__42191\
        );

    \I__9455\ : InMux
    port map (
            O => \N__42222\,
            I => \N__42191\
        );

    \I__9454\ : InMux
    port map (
            O => \N__42221\,
            I => \N__42191\
        );

    \I__9453\ : InMux
    port map (
            O => \N__42220\,
            I => \N__42191\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__42217\,
            I => \N__42186\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__42212\,
            I => \N__42186\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__42209\,
            I => \N__42183\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__42206\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__42203\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42200\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__42191\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__9445\ : Odrv4
    port map (
            O => \N__42186\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__9444\ : Odrv4
    port map (
            O => \N__42183\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__9443\ : InMux
    port map (
            O => \N__42170\,
            I => \N__42166\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42161\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__42166\,
            I => \N__42158\
        );

    \I__9440\ : CascadeMux
    port map (
            O => \N__42165\,
            I => \N__42155\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42164\,
            I => \N__42151\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__42161\,
            I => \N__42148\
        );

    \I__9437\ : Span4Mux_v
    port map (
            O => \N__42158\,
            I => \N__42145\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42155\,
            I => \N__42142\
        );

    \I__9435\ : InMux
    port map (
            O => \N__42154\,
            I => \N__42139\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__42151\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__9433\ : Odrv12
    port map (
            O => \N__42148\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__42145\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__42142\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__42139\,
            I => \elapsed_time_ns_1_RNIRHL2M1_0_3\
        );

    \I__9429\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42125\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__42125\,
            I => \N__42122\
        );

    \I__9427\ : Odrv4
    port map (
            O => \N__42122\,
            I => \phase_controller_inst2.stoper_tr.un6_running_3\
        );

    \I__9426\ : CEMux
    port map (
            O => \N__42119\,
            I => \N__42112\
        );

    \I__9425\ : CEMux
    port map (
            O => \N__42118\,
            I => \N__42109\
        );

    \I__9424\ : CEMux
    port map (
            O => \N__42117\,
            I => \N__42106\
        );

    \I__9423\ : CEMux
    port map (
            O => \N__42116\,
            I => \N__42103\
        );

    \I__9422\ : CEMux
    port map (
            O => \N__42115\,
            I => \N__42099\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__42112\,
            I => \N__42084\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__42109\,
            I => \N__42076\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__42106\,
            I => \N__42076\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__42103\,
            I => \N__42073\
        );

    \I__9417\ : InMux
    port map (
            O => \N__42102\,
            I => \N__42066\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__42099\,
            I => \N__42063\
        );

    \I__9415\ : CEMux
    port map (
            O => \N__42098\,
            I => \N__42060\
        );

    \I__9414\ : InMux
    port map (
            O => \N__42097\,
            I => \N__42051\
        );

    \I__9413\ : InMux
    port map (
            O => \N__42096\,
            I => \N__42051\
        );

    \I__9412\ : InMux
    port map (
            O => \N__42095\,
            I => \N__42051\
        );

    \I__9411\ : InMux
    port map (
            O => \N__42094\,
            I => \N__42051\
        );

    \I__9410\ : InMux
    port map (
            O => \N__42093\,
            I => \N__42048\
        );

    \I__9409\ : InMux
    port map (
            O => \N__42092\,
            I => \N__42039\
        );

    \I__9408\ : InMux
    port map (
            O => \N__42091\,
            I => \N__42039\
        );

    \I__9407\ : InMux
    port map (
            O => \N__42090\,
            I => \N__42039\
        );

    \I__9406\ : InMux
    port map (
            O => \N__42089\,
            I => \N__42039\
        );

    \I__9405\ : InMux
    port map (
            O => \N__42088\,
            I => \N__42034\
        );

    \I__9404\ : InMux
    port map (
            O => \N__42087\,
            I => \N__42034\
        );

    \I__9403\ : Span4Mux_v
    port map (
            O => \N__42084\,
            I => \N__42031\
        );

    \I__9402\ : InMux
    port map (
            O => \N__42083\,
            I => \N__42024\
        );

    \I__9401\ : InMux
    port map (
            O => \N__42082\,
            I => \N__42024\
        );

    \I__9400\ : InMux
    port map (
            O => \N__42081\,
            I => \N__42024\
        );

    \I__9399\ : Span4Mux_v
    port map (
            O => \N__42076\,
            I => \N__42019\
        );

    \I__9398\ : Span4Mux_v
    port map (
            O => \N__42073\,
            I => \N__42019\
        );

    \I__9397\ : InMux
    port map (
            O => \N__42072\,
            I => \N__42010\
        );

    \I__9396\ : InMux
    port map (
            O => \N__42071\,
            I => \N__42010\
        );

    \I__9395\ : InMux
    port map (
            O => \N__42070\,
            I => \N__42010\
        );

    \I__9394\ : InMux
    port map (
            O => \N__42069\,
            I => \N__42010\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__42066\,
            I => \N__42007\
        );

    \I__9392\ : Span4Mux_v
    port map (
            O => \N__42063\,
            I => \N__42004\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__42060\,
            I => \N__42001\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__42051\,
            I => \N__41994\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__42048\,
            I => \N__41994\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__42039\,
            I => \N__41994\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__42034\,
            I => \N__41991\
        );

    \I__9386\ : Span4Mux_h
    port map (
            O => \N__42031\,
            I => \N__41982\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__42024\,
            I => \N__41982\
        );

    \I__9384\ : Span4Mux_v
    port map (
            O => \N__42019\,
            I => \N__41982\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__42010\,
            I => \N__41982\
        );

    \I__9382\ : Span4Mux_v
    port map (
            O => \N__42007\,
            I => \N__41979\
        );

    \I__9381\ : Span4Mux_v
    port map (
            O => \N__42004\,
            I => \N__41976\
        );

    \I__9380\ : Span12Mux_h
    port map (
            O => \N__42001\,
            I => \N__41973\
        );

    \I__9379\ : Span4Mux_v
    port map (
            O => \N__41994\,
            I => \N__41968\
        );

    \I__9378\ : Span4Mux_v
    port map (
            O => \N__41991\,
            I => \N__41968\
        );

    \I__9377\ : Span4Mux_h
    port map (
            O => \N__41982\,
            I => \N__41965\
        );

    \I__9376\ : Sp12to4
    port map (
            O => \N__41979\,
            I => \N__41960\
        );

    \I__9375\ : Sp12to4
    port map (
            O => \N__41976\,
            I => \N__41960\
        );

    \I__9374\ : Odrv12
    port map (
            O => \N__41973\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__9373\ : Odrv4
    port map (
            O => \N__41968\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__9372\ : Odrv4
    port map (
            O => \N__41965\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__9371\ : Odrv12
    port map (
            O => \N__41960\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__9370\ : InMux
    port map (
            O => \N__41951\,
            I => \N__41948\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__41948\,
            I => \N__41945\
        );

    \I__9368\ : Odrv4
    port map (
            O => \N__41945\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__9367\ : InMux
    port map (
            O => \N__41942\,
            I => \N__41939\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__41939\,
            I => \N__41936\
        );

    \I__9365\ : Odrv12
    port map (
            O => \N__41936\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41933\,
            I => \N__41930\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__41930\,
            I => \N__41927\
        );

    \I__9362\ : Odrv12
    port map (
            O => \N__41927\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__9361\ : InMux
    port map (
            O => \N__41924\,
            I => \N__41921\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__41921\,
            I => \N__41918\
        );

    \I__9359\ : Odrv12
    port map (
            O => \N__41918\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__9358\ : InMux
    port map (
            O => \N__41915\,
            I => \N__41912\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__41912\,
            I => \N__41909\
        );

    \I__9356\ : Odrv12
    port map (
            O => \N__41909\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__9355\ : CascadeMux
    port map (
            O => \N__41906\,
            I => \N__41903\
        );

    \I__9354\ : InMux
    port map (
            O => \N__41903\,
            I => \N__41900\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__41900\,
            I => \N__41897\
        );

    \I__9352\ : Span4Mux_v
    port map (
            O => \N__41897\,
            I => \N__41893\
        );

    \I__9351\ : InMux
    port map (
            O => \N__41896\,
            I => \N__41890\
        );

    \I__9350\ : Odrv4
    port map (
            O => \N__41893\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__41890\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__9348\ : InMux
    port map (
            O => \N__41885\,
            I => \N__41882\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__41882\,
            I => \N__41879\
        );

    \I__9346\ : Span4Mux_v
    port map (
            O => \N__41879\,
            I => \N__41874\
        );

    \I__9345\ : InMux
    port map (
            O => \N__41878\,
            I => \N__41869\
        );

    \I__9344\ : InMux
    port map (
            O => \N__41877\,
            I => \N__41869\
        );

    \I__9343\ : Span4Mux_h
    port map (
            O => \N__41874\,
            I => \N__41864\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__41869\,
            I => \N__41864\
        );

    \I__9341\ : Odrv4
    port map (
            O => \N__41864\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__9340\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41857\
        );

    \I__9339\ : InMux
    port map (
            O => \N__41860\,
            I => \N__41853\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__41857\,
            I => \N__41850\
        );

    \I__9337\ : InMux
    port map (
            O => \N__41856\,
            I => \N__41847\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__41853\,
            I => \N__41842\
        );

    \I__9335\ : Span4Mux_v
    port map (
            O => \N__41850\,
            I => \N__41837\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__41847\,
            I => \N__41837\
        );

    \I__9333\ : InMux
    port map (
            O => \N__41846\,
            I => \N__41832\
        );

    \I__9332\ : InMux
    port map (
            O => \N__41845\,
            I => \N__41832\
        );

    \I__9331\ : Odrv4
    port map (
            O => \N__41842\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__9330\ : Odrv4
    port map (
            O => \N__41837\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__41832\,
            I => \elapsed_time_ns_1_RNIFG4DM1_0_16\
        );

    \I__9328\ : CascadeMux
    port map (
            O => \N__41825\,
            I => \N__41817\
        );

    \I__9327\ : CascadeMux
    port map (
            O => \N__41824\,
            I => \N__41812\
        );

    \I__9326\ : CascadeMux
    port map (
            O => \N__41823\,
            I => \N__41806\
        );

    \I__9325\ : CascadeMux
    port map (
            O => \N__41822\,
            I => \N__41800\
        );

    \I__9324\ : CascadeMux
    port map (
            O => \N__41821\,
            I => \N__41797\
        );

    \I__9323\ : InMux
    port map (
            O => \N__41820\,
            I => \N__41793\
        );

    \I__9322\ : InMux
    port map (
            O => \N__41817\,
            I => \N__41790\
        );

    \I__9321\ : CascadeMux
    port map (
            O => \N__41816\,
            I => \N__41787\
        );

    \I__9320\ : CascadeMux
    port map (
            O => \N__41815\,
            I => \N__41783\
        );

    \I__9319\ : InMux
    port map (
            O => \N__41812\,
            I => \N__41780\
        );

    \I__9318\ : CascadeMux
    port map (
            O => \N__41811\,
            I => \N__41777\
        );

    \I__9317\ : CascadeMux
    port map (
            O => \N__41810\,
            I => \N__41774\
        );

    \I__9316\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41771\
        );

    \I__9315\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41765\
        );

    \I__9314\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41762\
        );

    \I__9313\ : InMux
    port map (
            O => \N__41804\,
            I => \N__41755\
        );

    \I__9312\ : InMux
    port map (
            O => \N__41803\,
            I => \N__41755\
        );

    \I__9311\ : InMux
    port map (
            O => \N__41800\,
            I => \N__41755\
        );

    \I__9310\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41747\
        );

    \I__9309\ : CascadeMux
    port map (
            O => \N__41796\,
            I => \N__41744\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__41793\,
            I => \N__41738\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__41790\,
            I => \N__41738\
        );

    \I__9306\ : InMux
    port map (
            O => \N__41787\,
            I => \N__41731\
        );

    \I__9305\ : InMux
    port map (
            O => \N__41786\,
            I => \N__41731\
        );

    \I__9304\ : InMux
    port map (
            O => \N__41783\,
            I => \N__41731\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__41780\,
            I => \N__41728\
        );

    \I__9302\ : InMux
    port map (
            O => \N__41777\,
            I => \N__41725\
        );

    \I__9301\ : InMux
    port map (
            O => \N__41774\,
            I => \N__41722\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__41771\,
            I => \N__41718\
        );

    \I__9299\ : CascadeMux
    port map (
            O => \N__41770\,
            I => \N__41715\
        );

    \I__9298\ : CascadeMux
    port map (
            O => \N__41769\,
            I => \N__41712\
        );

    \I__9297\ : CascadeMux
    port map (
            O => \N__41768\,
            I => \N__41709\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__41765\,
            I => \N__41706\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__41762\,
            I => \N__41701\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__41755\,
            I => \N__41701\
        );

    \I__9293\ : CascadeMux
    port map (
            O => \N__41754\,
            I => \N__41697\
        );

    \I__9292\ : CascadeMux
    port map (
            O => \N__41753\,
            I => \N__41694\
        );

    \I__9291\ : CascadeMux
    port map (
            O => \N__41752\,
            I => \N__41691\
        );

    \I__9290\ : CascadeMux
    port map (
            O => \N__41751\,
            I => \N__41686\
        );

    \I__9289\ : CascadeMux
    port map (
            O => \N__41750\,
            I => \N__41682\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__41747\,
            I => \N__41679\
        );

    \I__9287\ : InMux
    port map (
            O => \N__41744\,
            I => \N__41674\
        );

    \I__9286\ : InMux
    port map (
            O => \N__41743\,
            I => \N__41674\
        );

    \I__9285\ : Span4Mux_v
    port map (
            O => \N__41738\,
            I => \N__41669\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__41731\,
            I => \N__41669\
        );

    \I__9283\ : Span4Mux_v
    port map (
            O => \N__41728\,
            I => \N__41662\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__41725\,
            I => \N__41662\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__41722\,
            I => \N__41662\
        );

    \I__9280\ : InMux
    port map (
            O => \N__41721\,
            I => \N__41659\
        );

    \I__9279\ : Span4Mux_v
    port map (
            O => \N__41718\,
            I => \N__41656\
        );

    \I__9278\ : InMux
    port map (
            O => \N__41715\,
            I => \N__41653\
        );

    \I__9277\ : InMux
    port map (
            O => \N__41712\,
            I => \N__41650\
        );

    \I__9276\ : InMux
    port map (
            O => \N__41709\,
            I => \N__41647\
        );

    \I__9275\ : Span4Mux_h
    port map (
            O => \N__41706\,
            I => \N__41642\
        );

    \I__9274\ : Span4Mux_h
    port map (
            O => \N__41701\,
            I => \N__41642\
        );

    \I__9273\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41635\
        );

    \I__9272\ : InMux
    port map (
            O => \N__41697\,
            I => \N__41635\
        );

    \I__9271\ : InMux
    port map (
            O => \N__41694\,
            I => \N__41635\
        );

    \I__9270\ : InMux
    port map (
            O => \N__41691\,
            I => \N__41622\
        );

    \I__9269\ : InMux
    port map (
            O => \N__41690\,
            I => \N__41622\
        );

    \I__9268\ : InMux
    port map (
            O => \N__41689\,
            I => \N__41622\
        );

    \I__9267\ : InMux
    port map (
            O => \N__41686\,
            I => \N__41622\
        );

    \I__9266\ : InMux
    port map (
            O => \N__41685\,
            I => \N__41622\
        );

    \I__9265\ : InMux
    port map (
            O => \N__41682\,
            I => \N__41622\
        );

    \I__9264\ : Span4Mux_v
    port map (
            O => \N__41679\,
            I => \N__41617\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__41674\,
            I => \N__41617\
        );

    \I__9262\ : Span4Mux_h
    port map (
            O => \N__41669\,
            I => \N__41612\
        );

    \I__9261\ : Span4Mux_h
    port map (
            O => \N__41662\,
            I => \N__41612\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__41659\,
            I => \N__41609\
        );

    \I__9259\ : Odrv4
    port map (
            O => \N__41656\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__41653\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__41650\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__41647\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9255\ : Odrv4
    port map (
            O => \N__41642\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__41635\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__41622\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9252\ : Odrv4
    port map (
            O => \N__41617\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9251\ : Odrv4
    port map (
            O => \N__41612\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9250\ : Odrv12
    port map (
            O => \N__41609\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__9249\ : InMux
    port map (
            O => \N__41588\,
            I => \N__41579\
        );

    \I__9248\ : InMux
    port map (
            O => \N__41587\,
            I => \N__41576\
        );

    \I__9247\ : InMux
    port map (
            O => \N__41586\,
            I => \N__41573\
        );

    \I__9246\ : InMux
    port map (
            O => \N__41585\,
            I => \N__41570\
        );

    \I__9245\ : InMux
    port map (
            O => \N__41584\,
            I => \N__41565\
        );

    \I__9244\ : InMux
    port map (
            O => \N__41583\,
            I => \N__41565\
        );

    \I__9243\ : InMux
    port map (
            O => \N__41582\,
            I => \N__41562\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__41579\,
            I => \N__41556\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__41576\,
            I => \N__41556\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__41573\,
            I => \N__41552\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__41570\,
            I => \N__41547\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__41565\,
            I => \N__41547\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__41562\,
            I => \N__41544\
        );

    \I__9236\ : InMux
    port map (
            O => \N__41561\,
            I => \N__41541\
        );

    \I__9235\ : Span4Mux_v
    port map (
            O => \N__41556\,
            I => \N__41538\
        );

    \I__9234\ : InMux
    port map (
            O => \N__41555\,
            I => \N__41535\
        );

    \I__9233\ : Span4Mux_v
    port map (
            O => \N__41552\,
            I => \N__41530\
        );

    \I__9232\ : Span4Mux_v
    port map (
            O => \N__41547\,
            I => \N__41530\
        );

    \I__9231\ : Span4Mux_v
    port map (
            O => \N__41544\,
            I => \N__41525\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__41541\,
            I => \N__41525\
        );

    \I__9229\ : Odrv4
    port map (
            O => \N__41538\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__41535\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__9227\ : Odrv4
    port map (
            O => \N__41530\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__9226\ : Odrv4
    port map (
            O => \N__41525\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9\
        );

    \I__9225\ : InMux
    port map (
            O => \N__41516\,
            I => \N__41513\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__41513\,
            I => \N__41510\
        );

    \I__9223\ : Span4Mux_v
    port map (
            O => \N__41510\,
            I => \N__41507\
        );

    \I__9222\ : Odrv4
    port map (
            O => \N__41507\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16\
        );

    \I__9221\ : InMux
    port map (
            O => \N__41504\,
            I => \N__41500\
        );

    \I__9220\ : InMux
    port map (
            O => \N__41503\,
            I => \N__41493\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__41500\,
            I => \N__41490\
        );

    \I__9218\ : InMux
    port map (
            O => \N__41499\,
            I => \N__41487\
        );

    \I__9217\ : InMux
    port map (
            O => \N__41498\,
            I => \N__41484\
        );

    \I__9216\ : CascadeMux
    port map (
            O => \N__41497\,
            I => \N__41481\
        );

    \I__9215\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41476\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__41493\,
            I => \N__41469\
        );

    \I__9213\ : Span4Mux_h
    port map (
            O => \N__41490\,
            I => \N__41469\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__41487\,
            I => \N__41469\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__41484\,
            I => \N__41466\
        );

    \I__9210\ : InMux
    port map (
            O => \N__41481\,
            I => \N__41461\
        );

    \I__9209\ : InMux
    port map (
            O => \N__41480\,
            I => \N__41461\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41479\,
            I => \N__41458\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__41476\,
            I => \N__41453\
        );

    \I__9206\ : Span4Mux_v
    port map (
            O => \N__41469\,
            I => \N__41453\
        );

    \I__9205\ : Span4Mux_h
    port map (
            O => \N__41466\,
            I => \N__41450\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__41461\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__41458\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__9202\ : Odrv4
    port map (
            O => \N__41453\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__9201\ : Odrv4
    port map (
            O => \N__41450\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__9200\ : InMux
    port map (
            O => \N__41441\,
            I => \N__41438\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__41438\,
            I => \N__41435\
        );

    \I__9198\ : Odrv4
    port map (
            O => \N__41435\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1\
        );

    \I__9197\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41427\
        );

    \I__9196\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41422\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41430\,
            I => \N__41422\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__41427\,
            I => \N__41419\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__41422\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1\
        );

    \I__9192\ : Odrv4
    port map (
            O => \N__41419\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1\
        );

    \I__9191\ : InMux
    port map (
            O => \N__41414\,
            I => \N__41410\
        );

    \I__9190\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41407\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__41410\,
            I => \phase_controller_inst1.stoper_tr.N_235\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__41407\,
            I => \phase_controller_inst1.stoper_tr.N_235\
        );

    \I__9187\ : CascadeMux
    port map (
            O => \N__41402\,
            I => \elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_\
        );

    \I__9186\ : InMux
    port map (
            O => \N__41399\,
            I => \N__41396\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__41396\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\
        );

    \I__9184\ : CascadeMux
    port map (
            O => \N__41393\,
            I => \N__41390\
        );

    \I__9183\ : InMux
    port map (
            O => \N__41390\,
            I => \N__41387\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__41387\,
            I => \phase_controller_inst1.stoper_tr.un6_running_1\
        );

    \I__9181\ : InMux
    port map (
            O => \N__41384\,
            I => \N__41381\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__41381\,
            I => \N__41378\
        );

    \I__9179\ : Odrv4
    port map (
            O => \N__41378\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__9178\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41372\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__41372\,
            I => \N__41369\
        );

    \I__9176\ : Odrv12
    port map (
            O => \N__41369\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__9175\ : InMux
    port map (
            O => \N__41366\,
            I => \N__41363\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41363\,
            I => \N__41360\
        );

    \I__9173\ : Odrv12
    port map (
            O => \N__41360\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__9172\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41354\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__41354\,
            I => \N__41351\
        );

    \I__9170\ : Span4Mux_v
    port map (
            O => \N__41351\,
            I => \N__41348\
        );

    \I__9169\ : Odrv4
    port map (
            O => \N__41348\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__9168\ : InMux
    port map (
            O => \N__41345\,
            I => \N__41342\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__41342\,
            I => \N__41339\
        );

    \I__9166\ : Span4Mux_h
    port map (
            O => \N__41339\,
            I => \N__41336\
        );

    \I__9165\ : Odrv4
    port map (
            O => \N__41336\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41333\,
            I => \N__41330\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__41330\,
            I => \N__41327\
        );

    \I__9162\ : Odrv4
    port map (
            O => \N__41327\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41324\,
            I => \N__41321\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__41321\,
            I => \N__41318\
        );

    \I__9159\ : Odrv12
    port map (
            O => \N__41318\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__9158\ : InMux
    port map (
            O => \N__41315\,
            I => \N__41312\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__41312\,
            I => \N__41309\
        );

    \I__9156\ : Odrv12
    port map (
            O => \N__41309\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__9155\ : InMux
    port map (
            O => \N__41306\,
            I => \N__41303\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41303\,
            I => \N__41300\
        );

    \I__9153\ : Odrv12
    port map (
            O => \N__41300\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__9152\ : InMux
    port map (
            O => \N__41297\,
            I => \N__41294\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__41294\,
            I => \N__41291\
        );

    \I__9150\ : Odrv4
    port map (
            O => \N__41291\,
            I => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\
        );

    \I__9149\ : CascadeMux
    port map (
            O => \N__41288\,
            I => \N__41285\
        );

    \I__9148\ : InMux
    port map (
            O => \N__41285\,
            I => \N__41281\
        );

    \I__9147\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41278\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__41281\,
            I => \N__41273\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__41278\,
            I => \N__41273\
        );

    \I__9144\ : Span4Mux_v
    port map (
            O => \N__41273\,
            I => \N__41269\
        );

    \I__9143\ : InMux
    port map (
            O => \N__41272\,
            I => \N__41266\
        );

    \I__9142\ : Odrv4
    port map (
            O => \N__41269\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__41266\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9140\ : CascadeMux
    port map (
            O => \N__41261\,
            I => \N__41258\
        );

    \I__9139\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41255\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__41255\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41252\,
            I => \N__41249\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41249\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__9135\ : CascadeMux
    port map (
            O => \N__41246\,
            I => \N__41243\
        );

    \I__9134\ : InMux
    port map (
            O => \N__41243\,
            I => \N__41240\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__41240\,
            I => \N__41237\
        );

    \I__9132\ : Odrv4
    port map (
            O => \N__41237\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__9131\ : CascadeMux
    port map (
            O => \N__41234\,
            I => \N__41231\
        );

    \I__9130\ : InMux
    port map (
            O => \N__41231\,
            I => \N__41228\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__41228\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__9128\ : InMux
    port map (
            O => \N__41225\,
            I => \N__41222\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__41222\,
            I => \N__41219\
        );

    \I__9126\ : Odrv4
    port map (
            O => \N__41219\,
            I => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\
        );

    \I__9125\ : CascadeMux
    port map (
            O => \N__41216\,
            I => \N__41212\
        );

    \I__9124\ : CascadeMux
    port map (
            O => \N__41215\,
            I => \N__41209\
        );

    \I__9123\ : InMux
    port map (
            O => \N__41212\,
            I => \N__41205\
        );

    \I__9122\ : InMux
    port map (
            O => \N__41209\,
            I => \N__41202\
        );

    \I__9121\ : InMux
    port map (
            O => \N__41208\,
            I => \N__41199\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__41205\,
            I => \N__41196\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__41202\,
            I => \N__41193\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__41199\,
            I => \N__41190\
        );

    \I__9117\ : Span4Mux_h
    port map (
            O => \N__41196\,
            I => \N__41185\
        );

    \I__9116\ : Span4Mux_v
    port map (
            O => \N__41193\,
            I => \N__41185\
        );

    \I__9115\ : Span4Mux_v
    port map (
            O => \N__41190\,
            I => \N__41182\
        );

    \I__9114\ : Odrv4
    port map (
            O => \N__41185\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__9113\ : Odrv4
    port map (
            O => \N__41182\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__9112\ : CascadeMux
    port map (
            O => \N__41177\,
            I => \N__41174\
        );

    \I__9111\ : InMux
    port map (
            O => \N__41174\,
            I => \N__41171\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__41171\,
            I => \N__41168\
        );

    \I__9109\ : Odrv4
    port map (
            O => \N__41168\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__9108\ : InMux
    port map (
            O => \N__41165\,
            I => \N__41162\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__41162\,
            I => \N__41159\
        );

    \I__9106\ : Odrv12
    port map (
            O => \N__41159\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__9105\ : InMux
    port map (
            O => \N__41156\,
            I => \N__41152\
        );

    \I__9104\ : InMux
    port map (
            O => \N__41155\,
            I => \N__41149\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__41152\,
            I => \N__41145\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__41149\,
            I => \N__41142\
        );

    \I__9101\ : InMux
    port map (
            O => \N__41148\,
            I => \N__41139\
        );

    \I__9100\ : Span4Mux_h
    port map (
            O => \N__41145\,
            I => \N__41136\
        );

    \I__9099\ : Odrv12
    port map (
            O => \N__41142\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__41139\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9097\ : Odrv4
    port map (
            O => \N__41136\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9096\ : CascadeMux
    port map (
            O => \N__41129\,
            I => \N__41126\
        );

    \I__9095\ : InMux
    port map (
            O => \N__41126\,
            I => \N__41123\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41123\,
            I => \N__41120\
        );

    \I__9093\ : Span4Mux_h
    port map (
            O => \N__41120\,
            I => \N__41117\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__41117\,
            I => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41114\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41111\,
            I => \N__41108\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__41108\,
            I => \N__41103\
        );

    \I__9088\ : InMux
    port map (
            O => \N__41107\,
            I => \N__41098\
        );

    \I__9087\ : InMux
    port map (
            O => \N__41106\,
            I => \N__41098\
        );

    \I__9086\ : Span4Mux_h
    port map (
            O => \N__41103\,
            I => \N__41095\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__41098\,
            I => \N__41092\
        );

    \I__9084\ : Odrv4
    port map (
            O => \N__41095\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9083\ : Odrv12
    port map (
            O => \N__41092\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9082\ : InMux
    port map (
            O => \N__41087\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__9081\ : InMux
    port map (
            O => \N__41084\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41081\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__9079\ : InMux
    port map (
            O => \N__41078\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__9078\ : InMux
    port map (
            O => \N__41075\,
            I => \N__41072\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__41072\,
            I => \N__41068\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41071\,
            I => \N__41065\
        );

    \I__9075\ : Span4Mux_v
    port map (
            O => \N__41068\,
            I => \N__41061\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__41065\,
            I => \N__41058\
        );

    \I__9073\ : InMux
    port map (
            O => \N__41064\,
            I => \N__41055\
        );

    \I__9072\ : Odrv4
    port map (
            O => \N__41061\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__41058\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__41055\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9069\ : CascadeMux
    port map (
            O => \N__41048\,
            I => \N__41045\
        );

    \I__9068\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41042\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__41042\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__9066\ : InMux
    port map (
            O => \N__41039\,
            I => \N__41036\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__41036\,
            I => \N__41033\
        );

    \I__9064\ : Span4Mux_h
    port map (
            O => \N__41033\,
            I => \N__41030\
        );

    \I__9063\ : Odrv4
    port map (
            O => \N__41030\,
            I => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41027\,
            I => \N__41024\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__41024\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__41021\,
            I => \N__41018\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41018\,
            I => \N__41015\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__41015\,
            I => \N__41012\
        );

    \I__9057\ : Odrv4
    port map (
            O => \N__41012\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__9056\ : InMux
    port map (
            O => \N__41009\,
            I => \bfn_17_17_0_\
        );

    \I__9055\ : InMux
    port map (
            O => \N__41006\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41003\,
            I => \N__40999\
        );

    \I__9053\ : CascadeMux
    port map (
            O => \N__41002\,
            I => \N__40996\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__40999\,
            I => \N__40992\
        );

    \I__9051\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40987\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40995\,
            I => \N__40987\
        );

    \I__9049\ : Span4Mux_h
    port map (
            O => \N__40992\,
            I => \N__40984\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__40987\,
            I => \N__40981\
        );

    \I__9047\ : Odrv4
    port map (
            O => \N__40984\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9046\ : Odrv12
    port map (
            O => \N__40981\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9045\ : InMux
    port map (
            O => \N__40976\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__9044\ : InMux
    port map (
            O => \N__40973\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__9043\ : CascadeMux
    port map (
            O => \N__40970\,
            I => \N__40966\
        );

    \I__9042\ : InMux
    port map (
            O => \N__40969\,
            I => \N__40960\
        );

    \I__9041\ : InMux
    port map (
            O => \N__40966\,
            I => \N__40960\
        );

    \I__9040\ : InMux
    port map (
            O => \N__40965\,
            I => \N__40957\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__40960\,
            I => \N__40952\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__40957\,
            I => \N__40952\
        );

    \I__9037\ : Span4Mux_h
    port map (
            O => \N__40952\,
            I => \N__40949\
        );

    \I__9036\ : Odrv4
    port map (
            O => \N__40949\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9035\ : InMux
    port map (
            O => \N__40946\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__9034\ : InMux
    port map (
            O => \N__40943\,
            I => \N__40938\
        );

    \I__9033\ : InMux
    port map (
            O => \N__40942\,
            I => \N__40935\
        );

    \I__9032\ : InMux
    port map (
            O => \N__40941\,
            I => \N__40932\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__40938\,
            I => \N__40929\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__40935\,
            I => \N__40926\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__40932\,
            I => \N__40921\
        );

    \I__9028\ : Span4Mux_h
    port map (
            O => \N__40929\,
            I => \N__40921\
        );

    \I__9027\ : Odrv4
    port map (
            O => \N__40926\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9026\ : Odrv4
    port map (
            O => \N__40921\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9025\ : InMux
    port map (
            O => \N__40916\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__9024\ : InMux
    port map (
            O => \N__40913\,
            I => \N__40906\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40912\,
            I => \N__40906\
        );

    \I__9022\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40903\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__40906\,
            I => \N__40900\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__40903\,
            I => \N__40897\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__40900\,
            I => \N__40894\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__40897\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__40894\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9016\ : InMux
    port map (
            O => \N__40889\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__9015\ : InMux
    port map (
            O => \N__40886\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__9014\ : InMux
    port map (
            O => \N__40883\,
            I => \bfn_17_18_0_\
        );

    \I__9013\ : CascadeMux
    port map (
            O => \N__40880\,
            I => \N__40876\
        );

    \I__9012\ : InMux
    port map (
            O => \N__40879\,
            I => \N__40872\
        );

    \I__9011\ : InMux
    port map (
            O => \N__40876\,
            I => \N__40867\
        );

    \I__9010\ : InMux
    port map (
            O => \N__40875\,
            I => \N__40867\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__40872\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__40867\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9007\ : InMux
    port map (
            O => \N__40862\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40859\,
            I => \bfn_17_16_0_\
        );

    \I__9005\ : InMux
    port map (
            O => \N__40856\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__9004\ : InMux
    port map (
            O => \N__40853\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__9003\ : InMux
    port map (
            O => \N__40850\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__9002\ : InMux
    port map (
            O => \N__40847\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40844\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__9000\ : InMux
    port map (
            O => \N__40841\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__8999\ : InMux
    port map (
            O => \N__40838\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__8998\ : InMux
    port map (
            O => \N__40835\,
            I => \N__40832\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__40832\,
            I => \N__40829\
        );

    \I__8996\ : Sp12to4
    port map (
            O => \N__40829\,
            I => \N__40823\
        );

    \I__8995\ : CascadeMux
    port map (
            O => \N__40828\,
            I => \N__40820\
        );

    \I__8994\ : InMux
    port map (
            O => \N__40827\,
            I => \N__40817\
        );

    \I__8993\ : InMux
    port map (
            O => \N__40826\,
            I => \N__40814\
        );

    \I__8992\ : Span12Mux_v
    port map (
            O => \N__40823\,
            I => \N__40811\
        );

    \I__8991\ : InMux
    port map (
            O => \N__40820\,
            I => \N__40808\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__40817\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__40814\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8988\ : Odrv12
    port map (
            O => \N__40811\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__40808\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__8986\ : InMux
    port map (
            O => \N__40799\,
            I => \N__40793\
        );

    \I__8985\ : InMux
    port map (
            O => \N__40798\,
            I => \N__40793\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__40793\,
            I => \N__40789\
        );

    \I__8983\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40786\
        );

    \I__8982\ : Odrv4
    port map (
            O => \N__40789\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__40786\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__8980\ : InMux
    port map (
            O => \N__40781\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__8979\ : InMux
    port map (
            O => \N__40778\,
            I => \N__40775\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__40775\,
            I => \N__40771\
        );

    \I__8977\ : InMux
    port map (
            O => \N__40774\,
            I => \N__40768\
        );

    \I__8976\ : Span4Mux_v
    port map (
            O => \N__40771\,
            I => \N__40763\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__40768\,
            I => \N__40763\
        );

    \I__8974\ : Span4Mux_h
    port map (
            O => \N__40763\,
            I => \N__40759\
        );

    \I__8973\ : InMux
    port map (
            O => \N__40762\,
            I => \N__40756\
        );

    \I__8972\ : Odrv4
    port map (
            O => \N__40759\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__40756\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__8970\ : InMux
    port map (
            O => \N__40751\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__8969\ : InMux
    port map (
            O => \N__40748\,
            I => \N__40745\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__40745\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__8967\ : InMux
    port map (
            O => \N__40742\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__8966\ : InMux
    port map (
            O => \N__40739\,
            I => \N__40736\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__40736\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__8964\ : InMux
    port map (
            O => \N__40733\,
            I => \N__40726\
        );

    \I__8963\ : InMux
    port map (
            O => \N__40732\,
            I => \N__40726\
        );

    \I__8962\ : InMux
    port map (
            O => \N__40731\,
            I => \N__40723\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__40726\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__40723\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__8959\ : InMux
    port map (
            O => \N__40718\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__8958\ : InMux
    port map (
            O => \N__40715\,
            I => \N__40708\
        );

    \I__8957\ : InMux
    port map (
            O => \N__40714\,
            I => \N__40708\
        );

    \I__8956\ : InMux
    port map (
            O => \N__40713\,
            I => \N__40705\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__40708\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__40705\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__8953\ : InMux
    port map (
            O => \N__40700\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__8952\ : InMux
    port map (
            O => \N__40697\,
            I => \N__40690\
        );

    \I__8951\ : InMux
    port map (
            O => \N__40696\,
            I => \N__40690\
        );

    \I__8950\ : InMux
    port map (
            O => \N__40695\,
            I => \N__40687\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__40690\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__40687\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__8947\ : InMux
    port map (
            O => \N__40682\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__8946\ : CascadeMux
    port map (
            O => \N__40679\,
            I => \N__40676\
        );

    \I__8945\ : InMux
    port map (
            O => \N__40676\,
            I => \N__40673\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__40673\,
            I => \N__40670\
        );

    \I__8943\ : Span4Mux_h
    port map (
            O => \N__40670\,
            I => \N__40667\
        );

    \I__8942\ : Odrv4
    port map (
            O => \N__40667\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__8941\ : CascadeMux
    port map (
            O => \N__40664\,
            I => \N__40661\
        );

    \I__8940\ : InMux
    port map (
            O => \N__40661\,
            I => \N__40658\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__40658\,
            I => \N__40655\
        );

    \I__8938\ : Span4Mux_v
    port map (
            O => \N__40655\,
            I => \N__40652\
        );

    \I__8937\ : Span4Mux_v
    port map (
            O => \N__40652\,
            I => \N__40649\
        );

    \I__8936\ : Odrv4
    port map (
            O => \N__40649\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__8935\ : InMux
    port map (
            O => \N__40646\,
            I => \N__40643\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__40643\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__8933\ : CascadeMux
    port map (
            O => \N__40640\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__8932\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40633\
        );

    \I__8931\ : CascadeMux
    port map (
            O => \N__40636\,
            I => \N__40630\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__40633\,
            I => \N__40627\
        );

    \I__8929\ : InMux
    port map (
            O => \N__40630\,
            I => \N__40624\
        );

    \I__8928\ : Sp12to4
    port map (
            O => \N__40627\,
            I => \N__40619\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__40624\,
            I => \N__40619\
        );

    \I__8926\ : Span12Mux_v
    port map (
            O => \N__40619\,
            I => \N__40616\
        );

    \I__8925\ : Odrv12
    port map (
            O => \N__40616\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__8924\ : CascadeMux
    port map (
            O => \N__40613\,
            I => \N__40609\
        );

    \I__8923\ : InMux
    port map (
            O => \N__40612\,
            I => \N__40606\
        );

    \I__8922\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40602\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__40606\,
            I => \N__40598\
        );

    \I__8920\ : InMux
    port map (
            O => \N__40605\,
            I => \N__40595\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__40602\,
            I => \N__40592\
        );

    \I__8918\ : InMux
    port map (
            O => \N__40601\,
            I => \N__40589\
        );

    \I__8917\ : Span4Mux_v
    port map (
            O => \N__40598\,
            I => \N__40586\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__40595\,
            I => \N__40583\
        );

    \I__8915\ : Span4Mux_h
    port map (
            O => \N__40592\,
            I => \N__40578\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__40589\,
            I => \N__40578\
        );

    \I__8913\ : Sp12to4
    port map (
            O => \N__40586\,
            I => \N__40575\
        );

    \I__8912\ : Span4Mux_v
    port map (
            O => \N__40583\,
            I => \N__40572\
        );

    \I__8911\ : Odrv4
    port map (
            O => \N__40578\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__8910\ : Odrv12
    port map (
            O => \N__40575\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__8909\ : Odrv4
    port map (
            O => \N__40572\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__8908\ : CascadeMux
    port map (
            O => \N__40565\,
            I => \N__40562\
        );

    \I__8907\ : InMux
    port map (
            O => \N__40562\,
            I => \N__40559\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__40559\,
            I => \N__40556\
        );

    \I__8905\ : Span4Mux_h
    port map (
            O => \N__40556\,
            I => \N__40553\
        );

    \I__8904\ : Span4Mux_h
    port map (
            O => \N__40553\,
            I => \N__40550\
        );

    \I__8903\ : Odrv4
    port map (
            O => \N__40550\,
            I => \current_shift_inst.PI_CTRL.integrator_i_30\
        );

    \I__8902\ : InMux
    port map (
            O => \N__40547\,
            I => \N__40543\
        );

    \I__8901\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40540\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__40543\,
            I => \N__40537\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__40540\,
            I => \N__40533\
        );

    \I__8898\ : Span4Mux_v
    port map (
            O => \N__40537\,
            I => \N__40530\
        );

    \I__8897\ : InMux
    port map (
            O => \N__40536\,
            I => \N__40527\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__40533\,
            I => \N__40524\
        );

    \I__8895\ : Span4Mux_h
    port map (
            O => \N__40530\,
            I => \N__40521\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__40527\,
            I => \N__40512\
        );

    \I__8893\ : Span4Mux_h
    port map (
            O => \N__40524\,
            I => \N__40512\
        );

    \I__8892\ : Span4Mux_h
    port map (
            O => \N__40521\,
            I => \N__40512\
        );

    \I__8891\ : InMux
    port map (
            O => \N__40520\,
            I => \N__40507\
        );

    \I__8890\ : InMux
    port map (
            O => \N__40519\,
            I => \N__40507\
        );

    \I__8889\ : Odrv4
    port map (
            O => \N__40512\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__40507\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__8887\ : InMux
    port map (
            O => \N__40502\,
            I => \N__40499\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__40499\,
            I => \N__40496\
        );

    \I__8885\ : Span4Mux_v
    port map (
            O => \N__40496\,
            I => \N__40493\
        );

    \I__8884\ : Span4Mux_h
    port map (
            O => \N__40493\,
            I => \N__40490\
        );

    \I__8883\ : Span4Mux_h
    port map (
            O => \N__40490\,
            I => \N__40487\
        );

    \I__8882\ : Odrv4
    port map (
            O => \N__40487\,
            I => \current_shift_inst.PI_CTRL.integrator_i_13\
        );

    \I__8881\ : InMux
    port map (
            O => \N__40484\,
            I => \N__40481\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__40481\,
            I => \N__40476\
        );

    \I__8879\ : InMux
    port map (
            O => \N__40480\,
            I => \N__40472\
        );

    \I__8878\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40469\
        );

    \I__8877\ : Span12Mux_v
    port map (
            O => \N__40476\,
            I => \N__40466\
        );

    \I__8876\ : InMux
    port map (
            O => \N__40475\,
            I => \N__40463\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__40472\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__40469\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__8873\ : Odrv12
    port map (
            O => \N__40466\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__40463\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40451\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__40451\,
            I => \N__40448\
        );

    \I__8869\ : Span4Mux_v
    port map (
            O => \N__40448\,
            I => \N__40445\
        );

    \I__8868\ : Odrv4
    port map (
            O => \N__40445\,
            I => \phase_controller_inst1.stoper_tr.un6_running_18\
        );

    \I__8867\ : CascadeMux
    port map (
            O => \N__40442\,
            I => \N__40439\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40439\,
            I => \N__40436\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__40436\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__8864\ : InMux
    port map (
            O => \N__40433\,
            I => \N__40430\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__40430\,
            I => \N__40427\
        );

    \I__8862\ : Span4Mux_v
    port map (
            O => \N__40427\,
            I => \N__40424\
        );

    \I__8861\ : Odrv4
    port map (
            O => \N__40424\,
            I => \phase_controller_inst1.stoper_tr.un6_running_19\
        );

    \I__8860\ : CascadeMux
    port map (
            O => \N__40421\,
            I => \N__40418\
        );

    \I__8859\ : InMux
    port map (
            O => \N__40418\,
            I => \N__40415\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__40415\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__8857\ : InMux
    port map (
            O => \N__40412\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_19\
        );

    \I__8856\ : InMux
    port map (
            O => \N__40409\,
            I => \N__40406\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__40406\,
            I => \N__40403\
        );

    \I__8854\ : Span12Mux_h
    port map (
            O => \N__40403\,
            I => \N__40400\
        );

    \I__8853\ : Odrv12
    port map (
            O => \N__40400\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__8852\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40394\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__40394\,
            I => \N__40391\
        );

    \I__8850\ : Span4Mux_v
    port map (
            O => \N__40391\,
            I => \N__40388\
        );

    \I__8849\ : Odrv4
    port map (
            O => \N__40388\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__8848\ : CascadeMux
    port map (
            O => \N__40385\,
            I => \N__40382\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40382\,
            I => \N__40379\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__40379\,
            I => \N__40376\
        );

    \I__8845\ : Span4Mux_v
    port map (
            O => \N__40376\,
            I => \N__40373\
        );

    \I__8844\ : Odrv4
    port map (
            O => \N__40373\,
            I => \phase_controller_inst1.stoper_tr.un6_running_10\
        );

    \I__8843\ : InMux
    port map (
            O => \N__40370\,
            I => \N__40367\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__40367\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__8841\ : InMux
    port map (
            O => \N__40364\,
            I => \N__40361\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40361\,
            I => \N__40358\
        );

    \I__8839\ : Span4Mux_h
    port map (
            O => \N__40358\,
            I => \N__40355\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__40355\,
            I => \phase_controller_inst1.stoper_tr.un6_running_11\
        );

    \I__8837\ : CascadeMux
    port map (
            O => \N__40352\,
            I => \N__40349\
        );

    \I__8836\ : InMux
    port map (
            O => \N__40349\,
            I => \N__40346\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__40346\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40343\,
            I => \N__40340\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__40340\,
            I => \N__40337\
        );

    \I__8832\ : Span4Mux_h
    port map (
            O => \N__40337\,
            I => \N__40334\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__40334\,
            I => \phase_controller_inst1.stoper_tr.un6_running_12\
        );

    \I__8830\ : CascadeMux
    port map (
            O => \N__40331\,
            I => \N__40328\
        );

    \I__8829\ : InMux
    port map (
            O => \N__40328\,
            I => \N__40325\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__40325\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40322\,
            I => \N__40319\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__40319\,
            I => \N__40316\
        );

    \I__8825\ : Span4Mux_h
    port map (
            O => \N__40316\,
            I => \N__40313\
        );

    \I__8824\ : Odrv4
    port map (
            O => \N__40313\,
            I => \phase_controller_inst1.stoper_tr.un6_running_13\
        );

    \I__8823\ : CascadeMux
    port map (
            O => \N__40310\,
            I => \N__40307\
        );

    \I__8822\ : InMux
    port map (
            O => \N__40307\,
            I => \N__40304\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40304\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__8820\ : CascadeMux
    port map (
            O => \N__40301\,
            I => \N__40298\
        );

    \I__8819\ : InMux
    port map (
            O => \N__40298\,
            I => \N__40295\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__40295\,
            I => \N__40292\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__40292\,
            I => \N__40289\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__40289\,
            I => \phase_controller_inst1.stoper_tr.un6_running_14\
        );

    \I__8815\ : InMux
    port map (
            O => \N__40286\,
            I => \N__40283\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__40283\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40280\,
            I => \N__40277\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__40277\,
            I => \phase_controller_inst1.stoper_tr.un6_running_15\
        );

    \I__8811\ : CascadeMux
    port map (
            O => \N__40274\,
            I => \N__40271\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40271\,
            I => \N__40268\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__40268\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__8808\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40262\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__40262\,
            I => \phase_controller_inst1.stoper_tr.un6_running_16\
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__40259\,
            I => \N__40256\
        );

    \I__8805\ : InMux
    port map (
            O => \N__40256\,
            I => \N__40253\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__40253\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__8803\ : InMux
    port map (
            O => \N__40250\,
            I => \N__40247\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__40247\,
            I => \N__40244\
        );

    \I__8801\ : Span4Mux_h
    port map (
            O => \N__40244\,
            I => \N__40241\
        );

    \I__8800\ : Odrv4
    port map (
            O => \N__40241\,
            I => \phase_controller_inst1.stoper_tr.un6_running_17\
        );

    \I__8799\ : CascadeMux
    port map (
            O => \N__40238\,
            I => \N__40235\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40235\,
            I => \N__40232\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__40232\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__8796\ : CascadeMux
    port map (
            O => \N__40229\,
            I => \N__40226\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40226\,
            I => \N__40223\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40223\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__8793\ : InMux
    port map (
            O => \N__40220\,
            I => \N__40217\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__40217\,
            I => \phase_controller_inst1.stoper_tr.un6_running_3\
        );

    \I__8791\ : CascadeMux
    port map (
            O => \N__40214\,
            I => \N__40211\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40211\,
            I => \N__40208\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__40208\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__8788\ : CascadeMux
    port map (
            O => \N__40205\,
            I => \N__40202\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40202\,
            I => \N__40199\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__40199\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40196\,
            I => \N__40193\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__40193\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40190\,
            I => \N__40187\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__40187\,
            I => \N__40184\
        );

    \I__8781\ : Odrv4
    port map (
            O => \N__40184\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__8780\ : CascadeMux
    port map (
            O => \N__40181\,
            I => \N__40178\
        );

    \I__8779\ : InMux
    port map (
            O => \N__40178\,
            I => \N__40175\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__40175\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__8777\ : InMux
    port map (
            O => \N__40172\,
            I => \N__40169\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__40169\,
            I => \N__40166\
        );

    \I__8775\ : Span4Mux_h
    port map (
            O => \N__40166\,
            I => \N__40163\
        );

    \I__8774\ : Odrv4
    port map (
            O => \N__40163\,
            I => \phase_controller_inst1.stoper_tr.un6_running_8\
        );

    \I__8773\ : CascadeMux
    port map (
            O => \N__40160\,
            I => \N__40157\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40157\,
            I => \N__40154\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__40154\,
            I => \N__40151\
        );

    \I__8770\ : Odrv4
    port map (
            O => \N__40151\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__8769\ : InMux
    port map (
            O => \N__40148\,
            I => \N__40145\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__40145\,
            I => \phase_controller_inst1.stoper_tr.un6_running_9\
        );

    \I__8767\ : CascadeMux
    port map (
            O => \N__40142\,
            I => \N__40139\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40139\,
            I => \N__40136\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__40136\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40133\,
            I => \N__40128\
        );

    \I__8763\ : InMux
    port map (
            O => \N__40132\,
            I => \N__40124\
        );

    \I__8762\ : InMux
    port map (
            O => \N__40131\,
            I => \N__40121\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__40128\,
            I => \N__40118\
        );

    \I__8760\ : InMux
    port map (
            O => \N__40127\,
            I => \N__40115\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__40124\,
            I => \N__40110\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__40121\,
            I => \N__40110\
        );

    \I__8757\ : Odrv12
    port map (
            O => \N__40118\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__40115\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__8755\ : Odrv4
    port map (
            O => \N__40110\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__8754\ : InMux
    port map (
            O => \N__40103\,
            I => \N__40100\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__40100\,
            I => \N__40097\
        );

    \I__8752\ : Span4Mux_v
    port map (
            O => \N__40097\,
            I => \N__40092\
        );

    \I__8751\ : InMux
    port map (
            O => \N__40096\,
            I => \N__40089\
        );

    \I__8750\ : InMux
    port map (
            O => \N__40095\,
            I => \N__40086\
        );

    \I__8749\ : Odrv4
    port map (
            O => \N__40092\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__40089\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__40086\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__8746\ : CascadeMux
    port map (
            O => \N__40079\,
            I => \N__40072\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40078\,
            I => \N__40069\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40077\,
            I => \N__40063\
        );

    \I__8743\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40063\
        );

    \I__8742\ : InMux
    port map (
            O => \N__40075\,
            I => \N__40060\
        );

    \I__8741\ : InMux
    port map (
            O => \N__40072\,
            I => \N__40053\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__40069\,
            I => \N__40049\
        );

    \I__8739\ : CascadeMux
    port map (
            O => \N__40068\,
            I => \N__40046\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__40063\,
            I => \N__40040\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__40060\,
            I => \N__40040\
        );

    \I__8736\ : InMux
    port map (
            O => \N__40059\,
            I => \N__40023\
        );

    \I__8735\ : InMux
    port map (
            O => \N__40058\,
            I => \N__40023\
        );

    \I__8734\ : InMux
    port map (
            O => \N__40057\,
            I => \N__40023\
        );

    \I__8733\ : InMux
    port map (
            O => \N__40056\,
            I => \N__40020\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__40053\,
            I => \N__40017\
        );

    \I__8731\ : InMux
    port map (
            O => \N__40052\,
            I => \N__40014\
        );

    \I__8730\ : Span4Mux_v
    port map (
            O => \N__40049\,
            I => \N__40011\
        );

    \I__8729\ : InMux
    port map (
            O => \N__40046\,
            I => \N__40008\
        );

    \I__8728\ : InMux
    port map (
            O => \N__40045\,
            I => \N__40005\
        );

    \I__8727\ : Span4Mux_h
    port map (
            O => \N__40040\,
            I => \N__40002\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40039\,
            I => \N__39995\
        );

    \I__8725\ : InMux
    port map (
            O => \N__40038\,
            I => \N__39995\
        );

    \I__8724\ : InMux
    port map (
            O => \N__40037\,
            I => \N__39995\
        );

    \I__8723\ : InMux
    port map (
            O => \N__40036\,
            I => \N__39980\
        );

    \I__8722\ : InMux
    port map (
            O => \N__40035\,
            I => \N__39980\
        );

    \I__8721\ : InMux
    port map (
            O => \N__40034\,
            I => \N__39980\
        );

    \I__8720\ : InMux
    port map (
            O => \N__40033\,
            I => \N__39980\
        );

    \I__8719\ : InMux
    port map (
            O => \N__40032\,
            I => \N__39980\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40031\,
            I => \N__39980\
        );

    \I__8717\ : InMux
    port map (
            O => \N__40030\,
            I => \N__39980\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__40023\,
            I => \N__39975\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__40020\,
            I => \N__39975\
        );

    \I__8714\ : Span4Mux_v
    port map (
            O => \N__40017\,
            I => \N__39970\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__40014\,
            I => \N__39970\
        );

    \I__8712\ : Odrv4
    port map (
            O => \N__40011\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__40008\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__40005\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8709\ : Odrv4
    port map (
            O => \N__40002\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__39995\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__39980\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8706\ : Odrv4
    port map (
            O => \N__39975\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8705\ : Odrv4
    port map (
            O => \N__39970\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8704\ : CascadeMux
    port map (
            O => \N__39953\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\
        );

    \I__8703\ : InMux
    port map (
            O => \N__39950\,
            I => \N__39947\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__39947\,
            I => \N__39943\
        );

    \I__8701\ : InMux
    port map (
            O => \N__39946\,
            I => \N__39940\
        );

    \I__8700\ : Span4Mux_v
    port map (
            O => \N__39943\,
            I => \N__39935\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__39940\,
            I => \N__39935\
        );

    \I__8698\ : Odrv4
    port map (
            O => \N__39935\,
            I => \phase_controller_inst1.stoper_tr.N_251\
        );

    \I__8697\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39929\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__39929\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\
        );

    \I__8695\ : InMux
    port map (
            O => \N__39926\,
            I => \N__39922\
        );

    \I__8694\ : CascadeMux
    port map (
            O => \N__39925\,
            I => \N__39919\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__39922\,
            I => \N__39913\
        );

    \I__8692\ : InMux
    port map (
            O => \N__39919\,
            I => \N__39908\
        );

    \I__8691\ : InMux
    port map (
            O => \N__39918\,
            I => \N__39908\
        );

    \I__8690\ : InMux
    port map (
            O => \N__39917\,
            I => \N__39903\
        );

    \I__8689\ : InMux
    port map (
            O => \N__39916\,
            I => \N__39903\
        );

    \I__8688\ : Odrv4
    port map (
            O => \N__39913\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__39908\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__39903\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9\
        );

    \I__8685\ : CascadeMux
    port map (
            O => \N__39896\,
            I => \N__39893\
        );

    \I__8684\ : InMux
    port map (
            O => \N__39893\,
            I => \N__39886\
        );

    \I__8683\ : InMux
    port map (
            O => \N__39892\,
            I => \N__39883\
        );

    \I__8682\ : InMux
    port map (
            O => \N__39891\,
            I => \N__39880\
        );

    \I__8681\ : InMux
    port map (
            O => \N__39890\,
            I => \N__39875\
        );

    \I__8680\ : InMux
    port map (
            O => \N__39889\,
            I => \N__39875\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__39886\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__39883\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__39880\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__39875\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14\
        );

    \I__8675\ : CascadeMux
    port map (
            O => \N__39866\,
            I => \elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_\
        );

    \I__8674\ : InMux
    port map (
            O => \N__39863\,
            I => \N__39858\
        );

    \I__8673\ : InMux
    port map (
            O => \N__39862\,
            I => \N__39855\
        );

    \I__8672\ : InMux
    port map (
            O => \N__39861\,
            I => \N__39852\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__39858\,
            I => \phase_controller_inst1.stoper_tr.N_244\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__39855\,
            I => \phase_controller_inst1.stoper_tr.N_244\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__39852\,
            I => \phase_controller_inst1.stoper_tr.N_244\
        );

    \I__8668\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39841\
        );

    \I__8667\ : InMux
    port map (
            O => \N__39844\,
            I => \N__39836\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__39841\,
            I => \N__39833\
        );

    \I__8665\ : InMux
    port map (
            O => \N__39840\,
            I => \N__39830\
        );

    \I__8664\ : InMux
    port map (
            O => \N__39839\,
            I => \N__39827\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__39836\,
            I => \N__39824\
        );

    \I__8662\ : Odrv12
    port map (
            O => \N__39833\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__39830\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__39827\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__8659\ : Odrv4
    port map (
            O => \N__39824\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__8658\ : CascadeMux
    port map (
            O => \N__39815\,
            I => \N__39812\
        );

    \I__8657\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39808\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__39811\,
            I => \N__39803\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__39808\,
            I => \N__39797\
        );

    \I__8654\ : InMux
    port map (
            O => \N__39807\,
            I => \N__39794\
        );

    \I__8653\ : InMux
    port map (
            O => \N__39806\,
            I => \N__39791\
        );

    \I__8652\ : InMux
    port map (
            O => \N__39803\,
            I => \N__39786\
        );

    \I__8651\ : InMux
    port map (
            O => \N__39802\,
            I => \N__39786\
        );

    \I__8650\ : InMux
    port map (
            O => \N__39801\,
            I => \N__39781\
        );

    \I__8649\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39781\
        );

    \I__8648\ : Odrv4
    port map (
            O => \N__39797\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__39794\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__39791\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__39786\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__39781\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__8643\ : CascadeMux
    port map (
            O => \N__39770\,
            I => \phase_controller_inst1.stoper_tr.N_211_cascade_\
        );

    \I__8642\ : CascadeMux
    port map (
            O => \N__39767\,
            I => \N__39749\
        );

    \I__8641\ : CascadeMux
    port map (
            O => \N__39766\,
            I => \N__39746\
        );

    \I__8640\ : CascadeMux
    port map (
            O => \N__39765\,
            I => \N__39739\
        );

    \I__8639\ : CascadeMux
    port map (
            O => \N__39764\,
            I => \N__39736\
        );

    \I__8638\ : InMux
    port map (
            O => \N__39763\,
            I => \N__39725\
        );

    \I__8637\ : InMux
    port map (
            O => \N__39762\,
            I => \N__39725\
        );

    \I__8636\ : InMux
    port map (
            O => \N__39761\,
            I => \N__39725\
        );

    \I__8635\ : InMux
    port map (
            O => \N__39760\,
            I => \N__39716\
        );

    \I__8634\ : InMux
    port map (
            O => \N__39759\,
            I => \N__39716\
        );

    \I__8633\ : InMux
    port map (
            O => \N__39758\,
            I => \N__39716\
        );

    \I__8632\ : InMux
    port map (
            O => \N__39757\,
            I => \N__39716\
        );

    \I__8631\ : CascadeMux
    port map (
            O => \N__39756\,
            I => \N__39710\
        );

    \I__8630\ : InMux
    port map (
            O => \N__39755\,
            I => \N__39707\
        );

    \I__8629\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39696\
        );

    \I__8628\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39696\
        );

    \I__8627\ : InMux
    port map (
            O => \N__39752\,
            I => \N__39696\
        );

    \I__8626\ : InMux
    port map (
            O => \N__39749\,
            I => \N__39696\
        );

    \I__8625\ : InMux
    port map (
            O => \N__39746\,
            I => \N__39696\
        );

    \I__8624\ : InMux
    port map (
            O => \N__39745\,
            I => \N__39689\
        );

    \I__8623\ : InMux
    port map (
            O => \N__39744\,
            I => \N__39689\
        );

    \I__8622\ : InMux
    port map (
            O => \N__39743\,
            I => \N__39689\
        );

    \I__8621\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39678\
        );

    \I__8620\ : InMux
    port map (
            O => \N__39739\,
            I => \N__39678\
        );

    \I__8619\ : InMux
    port map (
            O => \N__39736\,
            I => \N__39678\
        );

    \I__8618\ : InMux
    port map (
            O => \N__39735\,
            I => \N__39678\
        );

    \I__8617\ : InMux
    port map (
            O => \N__39734\,
            I => \N__39678\
        );

    \I__8616\ : InMux
    port map (
            O => \N__39733\,
            I => \N__39673\
        );

    \I__8615\ : InMux
    port map (
            O => \N__39732\,
            I => \N__39673\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__39725\,
            I => \N__39670\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__39716\,
            I => \N__39667\
        );

    \I__8612\ : InMux
    port map (
            O => \N__39715\,
            I => \N__39664\
        );

    \I__8611\ : InMux
    port map (
            O => \N__39714\,
            I => \N__39659\
        );

    \I__8610\ : InMux
    port map (
            O => \N__39713\,
            I => \N__39659\
        );

    \I__8609\ : InMux
    port map (
            O => \N__39710\,
            I => \N__39656\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__39707\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__39696\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__39689\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__39678\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__39673\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8603\ : Odrv4
    port map (
            O => \N__39670\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8602\ : Odrv4
    port map (
            O => \N__39667\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__39664\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__39659\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__39656\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8598\ : CascadeMux
    port map (
            O => \N__39635\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6_cascade_\
        );

    \I__8597\ : CascadeMux
    port map (
            O => \N__39632\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_\
        );

    \I__8596\ : InMux
    port map (
            O => \N__39629\,
            I => \N__39626\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__39626\,
            I => \N__39623\
        );

    \I__8594\ : Span4Mux_h
    port map (
            O => \N__39623\,
            I => \N__39620\
        );

    \I__8593\ : Odrv4
    port map (
            O => \N__39620\,
            I => \phase_controller_inst2.stoper_tr.un6_running_1\
        );

    \I__8592\ : InMux
    port map (
            O => \N__39617\,
            I => \N__39614\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__39614\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__8590\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39608\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__39608\,
            I => \N__39605\
        );

    \I__8588\ : Span4Mux_h
    port map (
            O => \N__39605\,
            I => \N__39602\
        );

    \I__8587\ : Odrv4
    port map (
            O => \N__39602\,
            I => \phase_controller_inst2.stoper_tr.un6_running_8\
        );

    \I__8586\ : InMux
    port map (
            O => \N__39599\,
            I => \N__39596\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__39596\,
            I => \N__39593\
        );

    \I__8584\ : Span4Mux_h
    port map (
            O => \N__39593\,
            I => \N__39590\
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__39590\,
            I => \phase_controller_inst2.stoper_tr.un6_running_2\
        );

    \I__8582\ : InMux
    port map (
            O => \N__39587\,
            I => \N__39584\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__39584\,
            I => \N__39581\
        );

    \I__8580\ : Span4Mux_h
    port map (
            O => \N__39581\,
            I => \N__39578\
        );

    \I__8579\ : Odrv4
    port map (
            O => \N__39578\,
            I => \phase_controller_inst1.stoper_tr.N_219\
        );

    \I__8578\ : InMux
    port map (
            O => \N__39575\,
            I => \N__39571\
        );

    \I__8577\ : InMux
    port map (
            O => \N__39574\,
            I => \N__39568\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__39571\,
            I => \N__39565\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__39568\,
            I => \N__39559\
        );

    \I__8574\ : Span12Mux_v
    port map (
            O => \N__39565\,
            I => \N__39559\
        );

    \I__8573\ : InMux
    port map (
            O => \N__39564\,
            I => \N__39556\
        );

    \I__8572\ : Odrv12
    port map (
            O => \N__39559\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__39556\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__8570\ : InMux
    port map (
            O => \N__39551\,
            I => \N__39546\
        );

    \I__8569\ : InMux
    port map (
            O => \N__39550\,
            I => \N__39541\
        );

    \I__8568\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39541\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__39546\,
            I => \N__39538\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__39541\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2\
        );

    \I__8565\ : Odrv4
    port map (
            O => \N__39538\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2\
        );

    \I__8564\ : InMux
    port map (
            O => \N__39533\,
            I => \N__39530\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__39530\,
            I => \N__39527\
        );

    \I__8562\ : Span4Mux_v
    port map (
            O => \N__39527\,
            I => \N__39524\
        );

    \I__8561\ : Odrv4
    port map (
            O => \N__39524\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6\
        );

    \I__8560\ : InMux
    port map (
            O => \N__39521\,
            I => \N__39517\
        );

    \I__8559\ : InMux
    port map (
            O => \N__39520\,
            I => \N__39514\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__39517\,
            I => \N__39510\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__39514\,
            I => \N__39506\
        );

    \I__8556\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39503\
        );

    \I__8555\ : Span4Mux_v
    port map (
            O => \N__39510\,
            I => \N__39500\
        );

    \I__8554\ : InMux
    port map (
            O => \N__39509\,
            I => \N__39497\
        );

    \I__8553\ : Span4Mux_h
    port map (
            O => \N__39506\,
            I => \N__39494\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__39503\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__39500\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__39497\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__8549\ : Odrv4
    port map (
            O => \N__39494\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__8548\ : CascadeMux
    port map (
            O => \N__39485\,
            I => \elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_\
        );

    \I__8547\ : CascadeMux
    port map (
            O => \N__39482\,
            I => \N__39479\
        );

    \I__8546\ : InMux
    port map (
            O => \N__39479\,
            I => \N__39474\
        );

    \I__8545\ : InMux
    port map (
            O => \N__39478\,
            I => \N__39471\
        );

    \I__8544\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39468\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__39474\,
            I => \phase_controller_inst1.stoper_tr.N_247\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__39471\,
            I => \phase_controller_inst1.stoper_tr.N_247\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__39468\,
            I => \phase_controller_inst1.stoper_tr.N_247\
        );

    \I__8540\ : CascadeMux
    port map (
            O => \N__39461\,
            I => \phase_controller_inst1.stoper_tr.N_247_cascade_\
        );

    \I__8539\ : CascadeMux
    port map (
            O => \N__39458\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_\
        );

    \I__8538\ : InMux
    port map (
            O => \N__39455\,
            I => \N__39452\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__39452\,
            I => \N__39449\
        );

    \I__8536\ : Span4Mux_v
    port map (
            O => \N__39449\,
            I => \N__39446\
        );

    \I__8535\ : Odrv4
    port map (
            O => \N__39446\,
            I => \phase_controller_inst2.stoper_tr.un6_running_6\
        );

    \I__8534\ : InMux
    port map (
            O => \N__39443\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__8533\ : InMux
    port map (
            O => \N__39440\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__8532\ : InMux
    port map (
            O => \N__39437\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39434\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__8530\ : InMux
    port map (
            O => \N__39431\,
            I => \N__39393\
        );

    \I__8529\ : InMux
    port map (
            O => \N__39430\,
            I => \N__39393\
        );

    \I__8528\ : InMux
    port map (
            O => \N__39429\,
            I => \N__39393\
        );

    \I__8527\ : InMux
    port map (
            O => \N__39428\,
            I => \N__39393\
        );

    \I__8526\ : InMux
    port map (
            O => \N__39427\,
            I => \N__39388\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39426\,
            I => \N__39388\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39425\,
            I => \N__39379\
        );

    \I__8523\ : InMux
    port map (
            O => \N__39424\,
            I => \N__39379\
        );

    \I__8522\ : InMux
    port map (
            O => \N__39423\,
            I => \N__39379\
        );

    \I__8521\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39379\
        );

    \I__8520\ : InMux
    port map (
            O => \N__39421\,
            I => \N__39370\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39420\,
            I => \N__39370\
        );

    \I__8518\ : InMux
    port map (
            O => \N__39419\,
            I => \N__39370\
        );

    \I__8517\ : InMux
    port map (
            O => \N__39418\,
            I => \N__39370\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39417\,
            I => \N__39361\
        );

    \I__8515\ : InMux
    port map (
            O => \N__39416\,
            I => \N__39361\
        );

    \I__8514\ : InMux
    port map (
            O => \N__39415\,
            I => \N__39361\
        );

    \I__8513\ : InMux
    port map (
            O => \N__39414\,
            I => \N__39361\
        );

    \I__8512\ : InMux
    port map (
            O => \N__39413\,
            I => \N__39352\
        );

    \I__8511\ : InMux
    port map (
            O => \N__39412\,
            I => \N__39352\
        );

    \I__8510\ : InMux
    port map (
            O => \N__39411\,
            I => \N__39352\
        );

    \I__8509\ : InMux
    port map (
            O => \N__39410\,
            I => \N__39352\
        );

    \I__8508\ : InMux
    port map (
            O => \N__39409\,
            I => \N__39343\
        );

    \I__8507\ : InMux
    port map (
            O => \N__39408\,
            I => \N__39343\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39343\
        );

    \I__8505\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39343\
        );

    \I__8504\ : InMux
    port map (
            O => \N__39405\,
            I => \N__39334\
        );

    \I__8503\ : InMux
    port map (
            O => \N__39404\,
            I => \N__39334\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39403\,
            I => \N__39334\
        );

    \I__8501\ : InMux
    port map (
            O => \N__39402\,
            I => \N__39334\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__39393\,
            I => \N__39321\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__39388\,
            I => \N__39321\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__39379\,
            I => \N__39321\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__39370\,
            I => \N__39321\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__39361\,
            I => \N__39321\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__39352\,
            I => \N__39321\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__39343\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__39334\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8492\ : Odrv12
    port map (
            O => \N__39321\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8491\ : InMux
    port map (
            O => \N__39314\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__8490\ : CEMux
    port map (
            O => \N__39311\,
            I => \N__39307\
        );

    \I__8489\ : CEMux
    port map (
            O => \N__39310\,
            I => \N__39304\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__39307\,
            I => \N__39299\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__39304\,
            I => \N__39296\
        );

    \I__8486\ : CEMux
    port map (
            O => \N__39303\,
            I => \N__39293\
        );

    \I__8485\ : CEMux
    port map (
            O => \N__39302\,
            I => \N__39290\
        );

    \I__8484\ : Span4Mux_v
    port map (
            O => \N__39299\,
            I => \N__39285\
        );

    \I__8483\ : Span4Mux_v
    port map (
            O => \N__39296\,
            I => \N__39285\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__39293\,
            I => \N__39280\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__39290\,
            I => \N__39280\
        );

    \I__8480\ : Odrv4
    port map (
            O => \N__39285\,
            I => \current_shift_inst.timer_s1.N_167_i\
        );

    \I__8479\ : Odrv4
    port map (
            O => \N__39280\,
            I => \current_shift_inst.timer_s1.N_167_i\
        );

    \I__8478\ : InMux
    port map (
            O => \N__39275\,
            I => \N__39272\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__39272\,
            I => \N__39266\
        );

    \I__8476\ : InMux
    port map (
            O => \N__39271\,
            I => \N__39263\
        );

    \I__8475\ : InMux
    port map (
            O => \N__39270\,
            I => \N__39258\
        );

    \I__8474\ : InMux
    port map (
            O => \N__39269\,
            I => \N__39258\
        );

    \I__8473\ : Odrv4
    port map (
            O => \N__39266\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__39263\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__39258\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39251\,
            I => \N__39248\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__39248\,
            I => \N__39245\
        );

    \I__8468\ : Span4Mux_h
    port map (
            O => \N__39245\,
            I => \N__39242\
        );

    \I__8467\ : Span4Mux_v
    port map (
            O => \N__39242\,
            I => \N__39239\
        );

    \I__8466\ : Odrv4
    port map (
            O => \N__39239\,
            I => \phase_controller_inst2.stoper_tr.un6_running_19\
        );

    \I__8465\ : InMux
    port map (
            O => \N__39236\,
            I => \N__39233\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__39233\,
            I => \N__39230\
        );

    \I__8463\ : Span4Mux_h
    port map (
            O => \N__39230\,
            I => \N__39227\
        );

    \I__8462\ : Span4Mux_v
    port map (
            O => \N__39227\,
            I => \N__39224\
        );

    \I__8461\ : Odrv4
    port map (
            O => \N__39224\,
            I => \phase_controller_inst2.stoper_tr.un6_running_16\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39218\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__39218\,
            I => \N__39215\
        );

    \I__8458\ : Span4Mux_v
    port map (
            O => \N__39215\,
            I => \N__39212\
        );

    \I__8457\ : Odrv4
    port map (
            O => \N__39212\,
            I => \phase_controller_inst2.stoper_tr.un6_running_15\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39209\,
            I => \N__39206\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__39206\,
            I => \N__39203\
        );

    \I__8454\ : Span4Mux_v
    port map (
            O => \N__39203\,
            I => \N__39200\
        );

    \I__8453\ : Odrv4
    port map (
            O => \N__39200\,
            I => \phase_controller_inst2.stoper_tr.un6_running_7\
        );

    \I__8452\ : InMux
    port map (
            O => \N__39197\,
            I => \bfn_16_23_0_\
        );

    \I__8451\ : InMux
    port map (
            O => \N__39194\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39191\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39188\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__8448\ : InMux
    port map (
            O => \N__39185\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__8447\ : InMux
    port map (
            O => \N__39182\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__8446\ : InMux
    port map (
            O => \N__39179\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__8445\ : InMux
    port map (
            O => \N__39176\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__8444\ : InMux
    port map (
            O => \N__39173\,
            I => \bfn_16_24_0_\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39170\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__8442\ : InMux
    port map (
            O => \N__39167\,
            I => \bfn_16_22_0_\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39164\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__8440\ : InMux
    port map (
            O => \N__39161\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__8439\ : InMux
    port map (
            O => \N__39158\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__8438\ : InMux
    port map (
            O => \N__39155\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__8437\ : InMux
    port map (
            O => \N__39152\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__8436\ : InMux
    port map (
            O => \N__39149\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__8435\ : InMux
    port map (
            O => \N__39146\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39143\,
            I => \N__39138\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39142\,
            I => \N__39135\
        );

    \I__8432\ : InMux
    port map (
            O => \N__39141\,
            I => \N__39132\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__39138\,
            I => \N__39127\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__39135\,
            I => \N__39127\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__39132\,
            I => \N__39121\
        );

    \I__8428\ : Sp12to4
    port map (
            O => \N__39127\,
            I => \N__39121\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39126\,
            I => \N__39118\
        );

    \I__8426\ : Span12Mux_v
    port map (
            O => \N__39121\,
            I => \N__39115\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__39118\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__8424\ : Odrv12
    port map (
            O => \N__39115\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__8423\ : InMux
    port map (
            O => \N__39110\,
            I => \N__39107\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__39107\,
            I => \N__39104\
        );

    \I__8421\ : Span4Mux_h
    port map (
            O => \N__39104\,
            I => \N__39101\
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__39101\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__8419\ : InMux
    port map (
            O => \N__39098\,
            I => \N__39095\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__39095\,
            I => \N__39092\
        );

    \I__8417\ : Odrv4
    port map (
            O => \N__39092\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__8416\ : InMux
    port map (
            O => \N__39089\,
            I => \bfn_16_21_0_\
        );

    \I__8415\ : InMux
    port map (
            O => \N__39086\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__8414\ : InMux
    port map (
            O => \N__39083\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39080\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39077\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__8411\ : InMux
    port map (
            O => \N__39074\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__8410\ : InMux
    port map (
            O => \N__39071\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39068\,
            I => \N__39052\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39067\,
            I => \N__39049\
        );

    \I__8407\ : CascadeMux
    port map (
            O => \N__39066\,
            I => \N__39044\
        );

    \I__8406\ : CascadeMux
    port map (
            O => \N__39065\,
            I => \N__39040\
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__39064\,
            I => \N__39036\
        );

    \I__8404\ : CascadeMux
    port map (
            O => \N__39063\,
            I => \N__39024\
        );

    \I__8403\ : CascadeMux
    port map (
            O => \N__39062\,
            I => \N__39020\
        );

    \I__8402\ : CascadeMux
    port map (
            O => \N__39061\,
            I => \N__39016\
        );

    \I__8401\ : CascadeMux
    port map (
            O => \N__39060\,
            I => \N__39012\
        );

    \I__8400\ : InMux
    port map (
            O => \N__39059\,
            I => \N__38998\
        );

    \I__8399\ : InMux
    port map (
            O => \N__39058\,
            I => \N__38998\
        );

    \I__8398\ : InMux
    port map (
            O => \N__39057\,
            I => \N__38998\
        );

    \I__8397\ : InMux
    port map (
            O => \N__39056\,
            I => \N__38998\
        );

    \I__8396\ : CascadeMux
    port map (
            O => \N__39055\,
            I => \N__38986\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__39052\,
            I => \N__38982\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__39049\,
            I => \N__38979\
        );

    \I__8393\ : InMux
    port map (
            O => \N__39048\,
            I => \N__38976\
        );

    \I__8392\ : InMux
    port map (
            O => \N__39047\,
            I => \N__38960\
        );

    \I__8391\ : InMux
    port map (
            O => \N__39044\,
            I => \N__38960\
        );

    \I__8390\ : InMux
    port map (
            O => \N__39043\,
            I => \N__38960\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39040\,
            I => \N__38960\
        );

    \I__8388\ : InMux
    port map (
            O => \N__39039\,
            I => \N__38960\
        );

    \I__8387\ : InMux
    port map (
            O => \N__39036\,
            I => \N__38960\
        );

    \I__8386\ : InMux
    port map (
            O => \N__39035\,
            I => \N__38960\
        );

    \I__8385\ : InMux
    port map (
            O => \N__39034\,
            I => \N__38951\
        );

    \I__8384\ : InMux
    port map (
            O => \N__39033\,
            I => \N__38951\
        );

    \I__8383\ : InMux
    port map (
            O => \N__39032\,
            I => \N__38951\
        );

    \I__8382\ : InMux
    port map (
            O => \N__39031\,
            I => \N__38951\
        );

    \I__8381\ : InMux
    port map (
            O => \N__39030\,
            I => \N__38942\
        );

    \I__8380\ : InMux
    port map (
            O => \N__39029\,
            I => \N__38942\
        );

    \I__8379\ : InMux
    port map (
            O => \N__39028\,
            I => \N__38942\
        );

    \I__8378\ : InMux
    port map (
            O => \N__39027\,
            I => \N__38942\
        );

    \I__8377\ : InMux
    port map (
            O => \N__39024\,
            I => \N__38925\
        );

    \I__8376\ : InMux
    port map (
            O => \N__39023\,
            I => \N__38925\
        );

    \I__8375\ : InMux
    port map (
            O => \N__39020\,
            I => \N__38925\
        );

    \I__8374\ : InMux
    port map (
            O => \N__39019\,
            I => \N__38925\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39016\,
            I => \N__38925\
        );

    \I__8372\ : InMux
    port map (
            O => \N__39015\,
            I => \N__38925\
        );

    \I__8371\ : InMux
    port map (
            O => \N__39012\,
            I => \N__38925\
        );

    \I__8370\ : InMux
    port map (
            O => \N__39011\,
            I => \N__38925\
        );

    \I__8369\ : InMux
    port map (
            O => \N__39010\,
            I => \N__38919\
        );

    \I__8368\ : InMux
    port map (
            O => \N__39009\,
            I => \N__38912\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39008\,
            I => \N__38912\
        );

    \I__8366\ : InMux
    port map (
            O => \N__39007\,
            I => \N__38912\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__38998\,
            I => \N__38909\
        );

    \I__8364\ : InMux
    port map (
            O => \N__38997\,
            I => \N__38906\
        );

    \I__8363\ : InMux
    port map (
            O => \N__38996\,
            I => \N__38899\
        );

    \I__8362\ : InMux
    port map (
            O => \N__38995\,
            I => \N__38899\
        );

    \I__8361\ : InMux
    port map (
            O => \N__38994\,
            I => \N__38899\
        );

    \I__8360\ : InMux
    port map (
            O => \N__38993\,
            I => \N__38890\
        );

    \I__8359\ : InMux
    port map (
            O => \N__38992\,
            I => \N__38890\
        );

    \I__8358\ : InMux
    port map (
            O => \N__38991\,
            I => \N__38890\
        );

    \I__8357\ : InMux
    port map (
            O => \N__38990\,
            I => \N__38890\
        );

    \I__8356\ : InMux
    port map (
            O => \N__38989\,
            I => \N__38883\
        );

    \I__8355\ : InMux
    port map (
            O => \N__38986\,
            I => \N__38883\
        );

    \I__8354\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38883\
        );

    \I__8353\ : Span4Mux_s1_h
    port map (
            O => \N__38982\,
            I => \N__38876\
        );

    \I__8352\ : Span4Mux_s1_v
    port map (
            O => \N__38979\,
            I => \N__38876\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__38976\,
            I => \N__38876\
        );

    \I__8350\ : InMux
    port map (
            O => \N__38975\,
            I => \N__38873\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__38960\,
            I => \N__38868\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__38951\,
            I => \N__38868\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__38942\,
            I => \N__38863\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__38925\,
            I => \N__38863\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__38924\,
            I => \N__38859\
        );

    \I__8344\ : CascadeMux
    port map (
            O => \N__38923\,
            I => \N__38855\
        );

    \I__8343\ : CascadeMux
    port map (
            O => \N__38922\,
            I => \N__38851\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__38919\,
            I => \N__38845\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__38912\,
            I => \N__38845\
        );

    \I__8340\ : Span4Mux_v
    port map (
            O => \N__38909\,
            I => \N__38840\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__38906\,
            I => \N__38840\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__38899\,
            I => \N__38835\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__38890\,
            I => \N__38835\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__38883\,
            I => \N__38832\
        );

    \I__8335\ : Sp12to4
    port map (
            O => \N__38876\,
            I => \N__38829\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__38873\,
            I => \N__38826\
        );

    \I__8333\ : Span4Mux_v
    port map (
            O => \N__38868\,
            I => \N__38821\
        );

    \I__8332\ : Span4Mux_v
    port map (
            O => \N__38863\,
            I => \N__38821\
        );

    \I__8331\ : InMux
    port map (
            O => \N__38862\,
            I => \N__38806\
        );

    \I__8330\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38806\
        );

    \I__8329\ : InMux
    port map (
            O => \N__38858\,
            I => \N__38806\
        );

    \I__8328\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38806\
        );

    \I__8327\ : InMux
    port map (
            O => \N__38854\,
            I => \N__38806\
        );

    \I__8326\ : InMux
    port map (
            O => \N__38851\,
            I => \N__38806\
        );

    \I__8325\ : InMux
    port map (
            O => \N__38850\,
            I => \N__38806\
        );

    \I__8324\ : Sp12to4
    port map (
            O => \N__38845\,
            I => \N__38803\
        );

    \I__8323\ : Sp12to4
    port map (
            O => \N__38840\,
            I => \N__38800\
        );

    \I__8322\ : Span12Mux_s9_h
    port map (
            O => \N__38835\,
            I => \N__38795\
        );

    \I__8321\ : Span12Mux_v
    port map (
            O => \N__38832\,
            I => \N__38790\
        );

    \I__8320\ : Span12Mux_s11_v
    port map (
            O => \N__38829\,
            I => \N__38790\
        );

    \I__8319\ : Span12Mux_s11_v
    port map (
            O => \N__38826\,
            I => \N__38783\
        );

    \I__8318\ : Sp12to4
    port map (
            O => \N__38821\,
            I => \N__38783\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__38806\,
            I => \N__38783\
        );

    \I__8316\ : Span12Mux_s10_v
    port map (
            O => \N__38803\,
            I => \N__38780\
        );

    \I__8315\ : Span12Mux_v
    port map (
            O => \N__38800\,
            I => \N__38777\
        );

    \I__8314\ : InMux
    port map (
            O => \N__38799\,
            I => \N__38772\
        );

    \I__8313\ : InMux
    port map (
            O => \N__38798\,
            I => \N__38772\
        );

    \I__8312\ : Span12Mux_v
    port map (
            O => \N__38795\,
            I => \N__38769\
        );

    \I__8311\ : Span12Mux_h
    port map (
            O => \N__38790\,
            I => \N__38764\
        );

    \I__8310\ : Span12Mux_h
    port map (
            O => \N__38783\,
            I => \N__38764\
        );

    \I__8309\ : Span12Mux_h
    port map (
            O => \N__38780\,
            I => \N__38757\
        );

    \I__8308\ : Span12Mux_h
    port map (
            O => \N__38777\,
            I => \N__38757\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__38772\,
            I => \N__38757\
        );

    \I__8306\ : Odrv12
    port map (
            O => \N__38769\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8305\ : Odrv12
    port map (
            O => \N__38764\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8304\ : Odrv12
    port map (
            O => \N__38757\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8303\ : InMux
    port map (
            O => \N__38750\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__8302\ : CascadeMux
    port map (
            O => \N__38747\,
            I => \N__38744\
        );

    \I__8301\ : InMux
    port map (
            O => \N__38744\,
            I => \N__38741\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__38741\,
            I => \N__38737\
        );

    \I__8299\ : InMux
    port map (
            O => \N__38740\,
            I => \N__38730\
        );

    \I__8298\ : Span4Mux_h
    port map (
            O => \N__38737\,
            I => \N__38720\
        );

    \I__8297\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38711\
        );

    \I__8296\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38711\
        );

    \I__8295\ : InMux
    port map (
            O => \N__38734\,
            I => \N__38711\
        );

    \I__8294\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38711\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__38730\,
            I => \N__38708\
        );

    \I__8292\ : InMux
    port map (
            O => \N__38729\,
            I => \N__38693\
        );

    \I__8291\ : InMux
    port map (
            O => \N__38728\,
            I => \N__38693\
        );

    \I__8290\ : InMux
    port map (
            O => \N__38727\,
            I => \N__38693\
        );

    \I__8289\ : InMux
    port map (
            O => \N__38726\,
            I => \N__38693\
        );

    \I__8288\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38693\
        );

    \I__8287\ : InMux
    port map (
            O => \N__38724\,
            I => \N__38693\
        );

    \I__8286\ : InMux
    port map (
            O => \N__38723\,
            I => \N__38693\
        );

    \I__8285\ : Odrv4
    port map (
            O => \N__38720\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__38711\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__8283\ : Odrv4
    port map (
            O => \N__38708\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__38693\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__8281\ : CascadeMux
    port map (
            O => \N__38684\,
            I => \N__38681\
        );

    \I__8280\ : InMux
    port map (
            O => \N__38681\,
            I => \N__38678\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__38678\,
            I => \N__38675\
        );

    \I__8278\ : Odrv4
    port map (
            O => \N__38675\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__8277\ : InMux
    port map (
            O => \N__38672\,
            I => \N__38669\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__38669\,
            I => \N__38666\
        );

    \I__8275\ : Span4Mux_v
    port map (
            O => \N__38666\,
            I => \N__38663\
        );

    \I__8274\ : Span4Mux_h
    port map (
            O => \N__38663\,
            I => \N__38660\
        );

    \I__8273\ : Odrv4
    port map (
            O => \N__38660\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__8272\ : InMux
    port map (
            O => \N__38657\,
            I => \N__38654\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__38654\,
            I => \N__38651\
        );

    \I__8270\ : Span4Mux_h
    port map (
            O => \N__38651\,
            I => \N__38648\
        );

    \I__8269\ : Odrv4
    port map (
            O => \N__38648\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__8268\ : CascadeMux
    port map (
            O => \N__38645\,
            I => \N__38642\
        );

    \I__8267\ : InMux
    port map (
            O => \N__38642\,
            I => \N__38639\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__38639\,
            I => \N__38636\
        );

    \I__8265\ : Odrv4
    port map (
            O => \N__38636\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__8264\ : InMux
    port map (
            O => \N__38633\,
            I => \N__38630\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__38630\,
            I => \N__38627\
        );

    \I__8262\ : Odrv4
    port map (
            O => \N__38627\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__8261\ : InMux
    port map (
            O => \N__38624\,
            I => \N__38621\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__38621\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__38618\,
            I => \N__38615\
        );

    \I__8258\ : InMux
    port map (
            O => \N__38615\,
            I => \N__38612\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__38612\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__8256\ : CascadeMux
    port map (
            O => \N__38609\,
            I => \N__38606\
        );

    \I__8255\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38603\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__38603\,
            I => \N__38600\
        );

    \I__8253\ : Odrv4
    port map (
            O => \N__38600\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__8252\ : CascadeMux
    port map (
            O => \N__38597\,
            I => \N__38594\
        );

    \I__8251\ : InMux
    port map (
            O => \N__38594\,
            I => \N__38591\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__38591\,
            I => \N__38588\
        );

    \I__8249\ : Span4Mux_h
    port map (
            O => \N__38588\,
            I => \N__38585\
        );

    \I__8248\ : Odrv4
    port map (
            O => \N__38585\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__8247\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38579\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__38579\,
            I => \N__38574\
        );

    \I__8245\ : InMux
    port map (
            O => \N__38578\,
            I => \N__38569\
        );

    \I__8244\ : InMux
    port map (
            O => \N__38577\,
            I => \N__38569\
        );

    \I__8243\ : Span4Mux_h
    port map (
            O => \N__38574\,
            I => \N__38566\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__38569\,
            I => \N__38563\
        );

    \I__8241\ : Odrv4
    port map (
            O => \N__38566\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__38563\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__8239\ : CascadeMux
    port map (
            O => \N__38558\,
            I => \N__38554\
        );

    \I__8238\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38551\
        );

    \I__8237\ : InMux
    port map (
            O => \N__38554\,
            I => \N__38548\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__38551\,
            I => \N__38545\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__38548\,
            I => \N__38542\
        );

    \I__8234\ : Span4Mux_h
    port map (
            O => \N__38545\,
            I => \N__38537\
        );

    \I__8233\ : Span4Mux_h
    port map (
            O => \N__38542\,
            I => \N__38537\
        );

    \I__8232\ : Span4Mux_h
    port map (
            O => \N__38537\,
            I => \N__38534\
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__38534\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__8230\ : InMux
    port map (
            O => \N__38531\,
            I => \N__38528\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__38528\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__8228\ : CascadeMux
    port map (
            O => \N__38525\,
            I => \N__38522\
        );

    \I__8227\ : InMux
    port map (
            O => \N__38522\,
            I => \N__38519\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__38519\,
            I => \N__38516\
        );

    \I__8225\ : Odrv4
    port map (
            O => \N__38516\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__8224\ : InMux
    port map (
            O => \N__38513\,
            I => \N__38510\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__38510\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__8222\ : CascadeMux
    port map (
            O => \N__38507\,
            I => \N__38504\
        );

    \I__8221\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38501\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__38501\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__8219\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38495\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__38495\,
            I => \N__38492\
        );

    \I__8217\ : Span4Mux_v
    port map (
            O => \N__38492\,
            I => \N__38489\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__38489\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__8215\ : InMux
    port map (
            O => \N__38486\,
            I => \N__38483\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__38483\,
            I => \N__38480\
        );

    \I__8213\ : Odrv12
    port map (
            O => \N__38480\,
            I => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__38477\,
            I => \N__38474\
        );

    \I__8211\ : InMux
    port map (
            O => \N__38474\,
            I => \N__38471\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__38471\,
            I => \N__38468\
        );

    \I__8209\ : Odrv4
    port map (
            O => \N__38468\,
            I => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__38465\,
            I => \N__38462\
        );

    \I__8207\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38459\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__38459\,
            I => \N__38456\
        );

    \I__8205\ : Span4Mux_v
    port map (
            O => \N__38456\,
            I => \N__38453\
        );

    \I__8204\ : Span4Mux_h
    port map (
            O => \N__38453\,
            I => \N__38450\
        );

    \I__8203\ : Odrv4
    port map (
            O => \N__38450\,
            I => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\
        );

    \I__8202\ : InMux
    port map (
            O => \N__38447\,
            I => \N__38444\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__38444\,
            I => \N__38441\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__38441\,
            I => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\
        );

    \I__8199\ : InMux
    port map (
            O => \N__38438\,
            I => \N__38435\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__38435\,
            I => \N__38432\
        );

    \I__8197\ : Span4Mux_v
    port map (
            O => \N__38432\,
            I => \N__38429\
        );

    \I__8196\ : Span4Mux_v
    port map (
            O => \N__38429\,
            I => \N__38424\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38428\,
            I => \N__38421\
        );

    \I__8194\ : CascadeMux
    port map (
            O => \N__38427\,
            I => \N__38418\
        );

    \I__8193\ : Span4Mux_v
    port map (
            O => \N__38424\,
            I => \N__38414\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__38421\,
            I => \N__38411\
        );

    \I__8191\ : InMux
    port map (
            O => \N__38418\,
            I => \N__38406\
        );

    \I__8190\ : InMux
    port map (
            O => \N__38417\,
            I => \N__38406\
        );

    \I__8189\ : Odrv4
    port map (
            O => \N__38414\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8188\ : Odrv4
    port map (
            O => \N__38411\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__38406\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8186\ : InMux
    port map (
            O => \N__38399\,
            I => \N__38396\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38396\,
            I => \N__38391\
        );

    \I__8184\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38388\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38394\,
            I => \N__38385\
        );

    \I__8182\ : Span4Mux_h
    port map (
            O => \N__38391\,
            I => \N__38378\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__38388\,
            I => \N__38378\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__38385\,
            I => \N__38378\
        );

    \I__8179\ : Span4Mux_v
    port map (
            O => \N__38378\,
            I => \N__38375\
        );

    \I__8178\ : Span4Mux_v
    port map (
            O => \N__38375\,
            I => \N__38372\
        );

    \I__8177\ : Odrv4
    port map (
            O => \N__38372\,
            I => \il_min_comp1_D2\
        );

    \I__8176\ : CascadeMux
    port map (
            O => \N__38369\,
            I => \N__38366\
        );

    \I__8175\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38360\
        );

    \I__8174\ : InMux
    port map (
            O => \N__38365\,
            I => \N__38360\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__38360\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38357\,
            I => \N__38354\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__38354\,
            I => \N__38350\
        );

    \I__8170\ : InMux
    port map (
            O => \N__38353\,
            I => \N__38347\
        );

    \I__8169\ : Sp12to4
    port map (
            O => \N__38350\,
            I => \N__38344\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__38347\,
            I => \N__38341\
        );

    \I__8167\ : Odrv12
    port map (
            O => \N__38344\,
            I => \phase_controller_inst1.N_56\
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__38341\,
            I => \phase_controller_inst1.N_56\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38327\
        );

    \I__8164\ : InMux
    port map (
            O => \N__38335\,
            I => \N__38327\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38334\,
            I => \N__38327\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__38327\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__8161\ : CascadeMux
    port map (
            O => \N__38324\,
            I => \N__38321\
        );

    \I__8160\ : InMux
    port map (
            O => \N__38321\,
            I => \N__38318\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38318\,
            I => \N__38315\
        );

    \I__8158\ : Span4Mux_h
    port map (
            O => \N__38315\,
            I => \N__38312\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__38312\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__8156\ : CascadeMux
    port map (
            O => \N__38309\,
            I => \N__38306\
        );

    \I__8155\ : InMux
    port map (
            O => \N__38306\,
            I => \N__38303\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38303\,
            I => \N__38300\
        );

    \I__8153\ : Odrv4
    port map (
            O => \N__38300\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__8152\ : InMux
    port map (
            O => \N__38297\,
            I => \N__38294\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__38294\,
            I => \N__38291\
        );

    \I__8150\ : Odrv4
    port map (
            O => \N__38291\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__8149\ : CascadeMux
    port map (
            O => \N__38288\,
            I => \N__38285\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38285\,
            I => \N__38282\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__38282\,
            I => \N__38279\
        );

    \I__8146\ : Span4Mux_h
    port map (
            O => \N__38279\,
            I => \N__38276\
        );

    \I__8145\ : Span4Mux_v
    port map (
            O => \N__38276\,
            I => \N__38273\
        );

    \I__8144\ : Odrv4
    port map (
            O => \N__38273\,
            I => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\
        );

    \I__8143\ : InMux
    port map (
            O => \N__38270\,
            I => \N__38267\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__38267\,
            I => \N__38264\
        );

    \I__8141\ : Span4Mux_v
    port map (
            O => \N__38264\,
            I => \N__38261\
        );

    \I__8140\ : Odrv4
    port map (
            O => \N__38261\,
            I => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\
        );

    \I__8139\ : InMux
    port map (
            O => \N__38258\,
            I => \N__38255\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38255\,
            I => \N__38252\
        );

    \I__8137\ : Span4Mux_h
    port map (
            O => \N__38252\,
            I => \N__38249\
        );

    \I__8136\ : Odrv4
    port map (
            O => \N__38249\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\
        );

    \I__8135\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38242\
        );

    \I__8134\ : InMux
    port map (
            O => \N__38245\,
            I => \N__38239\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__38242\,
            I => \N__38234\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__38239\,
            I => \N__38231\
        );

    \I__8131\ : InMux
    port map (
            O => \N__38238\,
            I => \N__38226\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38237\,
            I => \N__38226\
        );

    \I__8129\ : Span4Mux_v
    port map (
            O => \N__38234\,
            I => \N__38221\
        );

    \I__8128\ : Span4Mux_v
    port map (
            O => \N__38231\,
            I => \N__38221\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__38226\,
            I => \N__38218\
        );

    \I__8126\ : Odrv4
    port map (
            O => \N__38221\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18\
        );

    \I__8125\ : Odrv12
    port map (
            O => \N__38218\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18\
        );

    \I__8124\ : CascadeMux
    port map (
            O => \N__38213\,
            I => \elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38210\,
            I => \N__38207\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__38207\,
            I => \phase_controller_inst2.stoper_tr.un6_running_18\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38200\
        );

    \I__8120\ : InMux
    port map (
            O => \N__38203\,
            I => \N__38197\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__38200\,
            I => \N__38190\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__38197\,
            I => \N__38190\
        );

    \I__8117\ : InMux
    port map (
            O => \N__38196\,
            I => \N__38185\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38195\,
            I => \N__38185\
        );

    \I__8115\ : Odrv12
    port map (
            O => \N__38190\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38185\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17\
        );

    \I__8113\ : InMux
    port map (
            O => \N__38180\,
            I => \N__38177\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__38177\,
            I => \phase_controller_inst2.stoper_tr.un6_running_17\
        );

    \I__8111\ : CascadeMux
    port map (
            O => \N__38174\,
            I => \N__38171\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38171\,
            I => \N__38164\
        );

    \I__8109\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38161\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38169\,
            I => \N__38158\
        );

    \I__8107\ : InMux
    port map (
            O => \N__38168\,
            I => \N__38153\
        );

    \I__8106\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38153\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__38164\,
            I => \N__38150\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__38161\,
            I => \N__38147\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__38158\,
            I => \N__38144\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__38153\,
            I => \N__38139\
        );

    \I__8101\ : Span4Mux_h
    port map (
            O => \N__38150\,
            I => \N__38139\
        );

    \I__8100\ : Span4Mux_v
    port map (
            O => \N__38147\,
            I => \N__38136\
        );

    \I__8099\ : Span4Mux_h
    port map (
            O => \N__38144\,
            I => \N__38131\
        );

    \I__8098\ : Span4Mux_v
    port map (
            O => \N__38139\,
            I => \N__38131\
        );

    \I__8097\ : Odrv4
    port map (
            O => \N__38136\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__8096\ : Odrv4
    port map (
            O => \N__38131\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__8095\ : InMux
    port map (
            O => \N__38126\,
            I => \N__38123\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__38123\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9\
        );

    \I__8093\ : CascadeMux
    port map (
            O => \N__38120\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\
        );

    \I__8092\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38114\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__38114\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\
        );

    \I__8090\ : InMux
    port map (
            O => \N__38111\,
            I => \N__38105\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38110\,
            I => \N__38102\
        );

    \I__8088\ : CascadeMux
    port map (
            O => \N__38109\,
            I => \N__38099\
        );

    \I__8087\ : CascadeMux
    port map (
            O => \N__38108\,
            I => \N__38096\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__38105\,
            I => \N__38084\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__38102\,
            I => \N__38084\
        );

    \I__8084\ : InMux
    port map (
            O => \N__38099\,
            I => \N__38079\
        );

    \I__8083\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38079\
        );

    \I__8082\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38068\
        );

    \I__8081\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38068\
        );

    \I__8080\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38068\
        );

    \I__8079\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38068\
        );

    \I__8078\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38068\
        );

    \I__8077\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38063\
        );

    \I__8076\ : InMux
    port map (
            O => \N__38089\,
            I => \N__38063\
        );

    \I__8075\ : Span4Mux_v
    port map (
            O => \N__38084\,
            I => \N__38060\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__38079\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__38068\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__38063\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__8071\ : Odrv4
    port map (
            O => \N__38060\,
            I => \phase_controller_inst1.stoper_tr.N_241\
        );

    \I__8070\ : CascadeMux
    port map (
            O => \N__38051\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\
        );

    \I__8069\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38045\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__38045\,
            I => \phase_controller_inst2.stoper_tr.un6_running_9\
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__38042\,
            I => \N__38039\
        );

    \I__8066\ : InMux
    port map (
            O => \N__38039\,
            I => \N__38036\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__38036\,
            I => \N__38033\
        );

    \I__8064\ : Span4Mux_v
    port map (
            O => \N__38033\,
            I => \N__38029\
        );

    \I__8063\ : InMux
    port map (
            O => \N__38032\,
            I => \N__38026\
        );

    \I__8062\ : Odrv4
    port map (
            O => \N__38029\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__38026\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__8060\ : InMux
    port map (
            O => \N__38021\,
            I => \N__38018\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__38018\,
            I => \N__38015\
        );

    \I__8058\ : Span4Mux_v
    port map (
            O => \N__38015\,
            I => \N__38011\
        );

    \I__8057\ : InMux
    port map (
            O => \N__38014\,
            I => \N__38008\
        );

    \I__8056\ : Odrv4
    port map (
            O => \N__38011\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__38008\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__8054\ : InMux
    port map (
            O => \N__38003\,
            I => \N__38000\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__38000\,
            I => \elapsed_time_ns_1_RNIRAIF91_0_21\
        );

    \I__8052\ : InMux
    port map (
            O => \N__37997\,
            I => \N__37993\
        );

    \I__8051\ : InMux
    port map (
            O => \N__37996\,
            I => \N__37990\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__37993\,
            I => \N__37987\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__37990\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__8048\ : Odrv4
    port map (
            O => \N__37987\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__8047\ : InMux
    port map (
            O => \N__37982\,
            I => \N__37978\
        );

    \I__8046\ : InMux
    port map (
            O => \N__37981\,
            I => \N__37975\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__37978\,
            I => \elapsed_time_ns_1_RNI3JIF91_0_29\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__37975\,
            I => \elapsed_time_ns_1_RNI3JIF91_0_29\
        );

    \I__8043\ : CascadeMux
    port map (
            O => \N__37970\,
            I => \elapsed_time_ns_1_RNIRAIF91_0_21_cascade_\
        );

    \I__8042\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37964\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__37964\,
            I => \N__37960\
        );

    \I__8040\ : InMux
    port map (
            O => \N__37963\,
            I => \N__37957\
        );

    \I__8039\ : Span4Mux_h
    port map (
            O => \N__37960\,
            I => \N__37954\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__37957\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20\
        );

    \I__8037\ : Odrv4
    port map (
            O => \N__37954\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20\
        );

    \I__8036\ : InMux
    port map (
            O => \N__37949\,
            I => \N__37943\
        );

    \I__8035\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37943\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__37943\,
            I => \elapsed_time_ns_1_RNISBIF91_0_22\
        );

    \I__8033\ : InMux
    port map (
            O => \N__37940\,
            I => \N__37937\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__37937\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15\
        );

    \I__8031\ : CascadeMux
    port map (
            O => \N__37934\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_\
        );

    \I__8030\ : InMux
    port map (
            O => \N__37931\,
            I => \N__37928\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__37928\,
            I => \N__37925\
        );

    \I__8028\ : Span4Mux_h
    port map (
            O => \N__37925\,
            I => \N__37922\
        );

    \I__8027\ : Odrv4
    port map (
            O => \N__37922\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\
        );

    \I__8026\ : CascadeMux
    port map (
            O => \N__37919\,
            I => \phase_controller_inst1.stoper_tr.N_241_cascade_\
        );

    \I__8025\ : InMux
    port map (
            O => \N__37916\,
            I => \N__37913\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__37913\,
            I => \N__37910\
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__37910\,
            I => \phase_controller_inst2.stoper_tr.un6_running_14\
        );

    \I__8022\ : CascadeMux
    port map (
            O => \N__37907\,
            I => \N__37904\
        );

    \I__8021\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37899\
        );

    \I__8020\ : CascadeMux
    port map (
            O => \N__37903\,
            I => \N__37896\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__37902\,
            I => \N__37893\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__37899\,
            I => \N__37890\
        );

    \I__8017\ : InMux
    port map (
            O => \N__37896\,
            I => \N__37884\
        );

    \I__8016\ : InMux
    port map (
            O => \N__37893\,
            I => \N__37884\
        );

    \I__8015\ : Span4Mux_v
    port map (
            O => \N__37890\,
            I => \N__37881\
        );

    \I__8014\ : InMux
    port map (
            O => \N__37889\,
            I => \N__37878\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__37884\,
            I => \N__37875\
        );

    \I__8012\ : Odrv4
    port map (
            O => \N__37881\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__37878\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__8010\ : Odrv4
    port map (
            O => \N__37875\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__8009\ : InMux
    port map (
            O => \N__37868\,
            I => \N__37865\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__37865\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14\
        );

    \I__8007\ : InMux
    port map (
            O => \N__37862\,
            I => \N__37859\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__37859\,
            I => \N__37856\
        );

    \I__8005\ : Span4Mux_h
    port map (
            O => \N__37856\,
            I => \N__37853\
        );

    \I__8004\ : Odrv4
    port map (
            O => \N__37853\,
            I => \phase_controller_inst2.stoper_tr.un6_running_10\
        );

    \I__8003\ : CascadeMux
    port map (
            O => \N__37850\,
            I => \N__37847\
        );

    \I__8002\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37844\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__37844\,
            I => \N__37841\
        );

    \I__8000\ : Odrv4
    port map (
            O => \N__37841\,
            I => \phase_controller_inst2.stoper_tr.un6_running_11\
        );

    \I__7999\ : CascadeMux
    port map (
            O => \N__37838\,
            I => \N__37835\
        );

    \I__7998\ : InMux
    port map (
            O => \N__37835\,
            I => \N__37832\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__37832\,
            I => \N__37829\
        );

    \I__7996\ : Odrv4
    port map (
            O => \N__37829\,
            I => \phase_controller_inst2.stoper_tr.un6_running_12\
        );

    \I__7995\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37823\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__37823\,
            I => \N__37820\
        );

    \I__7993\ : Odrv4
    port map (
            O => \N__37820\,
            I => \phase_controller_inst2.stoper_tr.un6_running_13\
        );

    \I__7992\ : InMux
    port map (
            O => \N__37817\,
            I => \N__37812\
        );

    \I__7991\ : InMux
    port map (
            O => \N__37816\,
            I => \N__37809\
        );

    \I__7990\ : InMux
    port map (
            O => \N__37815\,
            I => \N__37806\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__37812\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__37809\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__37806\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__7986\ : CascadeMux
    port map (
            O => \N__37799\,
            I => \N__37794\
        );

    \I__7985\ : InMux
    port map (
            O => \N__37798\,
            I => \N__37790\
        );

    \I__7984\ : InMux
    port map (
            O => \N__37797\,
            I => \N__37787\
        );

    \I__7983\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37784\
        );

    \I__7982\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37781\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__37790\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__37787\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__37784\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__37781\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__7977\ : CascadeMux
    port map (
            O => \N__37772\,
            I => \N__37766\
        );

    \I__7976\ : InMux
    port map (
            O => \N__37771\,
            I => \N__37763\
        );

    \I__7975\ : InMux
    port map (
            O => \N__37770\,
            I => \N__37760\
        );

    \I__7974\ : InMux
    port map (
            O => \N__37769\,
            I => \N__37757\
        );

    \I__7973\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37754\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__37763\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__37760\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__37757\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__37754\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__7968\ : InMux
    port map (
            O => \N__37745\,
            I => \N__37739\
        );

    \I__7967\ : InMux
    port map (
            O => \N__37744\,
            I => \N__37736\
        );

    \I__7966\ : InMux
    port map (
            O => \N__37743\,
            I => \N__37733\
        );

    \I__7965\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37730\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__37739\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__37736\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__37733\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__37730\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__7960\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37717\
        );

    \I__7959\ : InMux
    port map (
            O => \N__37720\,
            I => \N__37713\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__37717\,
            I => \N__37710\
        );

    \I__7957\ : InMux
    port map (
            O => \N__37716\,
            I => \N__37707\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__37713\,
            I => \N__37704\
        );

    \I__7955\ : Odrv4
    port map (
            O => \N__37710\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__37707\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__37704\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__7952\ : CascadeMux
    port map (
            O => \N__37697\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\
        );

    \I__7951\ : CascadeMux
    port map (
            O => \N__37694\,
            I => \N__37691\
        );

    \I__7950\ : InMux
    port map (
            O => \N__37691\,
            I => \N__37688\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__37688\,
            I => \N__37683\
        );

    \I__7948\ : InMux
    port map (
            O => \N__37687\,
            I => \N__37678\
        );

    \I__7947\ : InMux
    port map (
            O => \N__37686\,
            I => \N__37678\
        );

    \I__7946\ : Span4Mux_h
    port map (
            O => \N__37683\,
            I => \N__37673\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__37678\,
            I => \N__37673\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__37673\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__7943\ : CascadeMux
    port map (
            O => \N__37670\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17_cascade_\
        );

    \I__7942\ : CascadeMux
    port map (
            O => \N__37667\,
            I => \elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_\
        );

    \I__7941\ : InMux
    port map (
            O => \N__37664\,
            I => \N__37661\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__37661\,
            I => \N__37658\
        );

    \I__7939\ : Span4Mux_h
    port map (
            O => \N__37658\,
            I => \N__37654\
        );

    \I__7938\ : InMux
    port map (
            O => \N__37657\,
            I => \N__37651\
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__37654\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__37651\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__7935\ : CascadeMux
    port map (
            O => \N__37646\,
            I => \elapsed_time_ns_1_RNICG2591_0_4_cascade_\
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__37643\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_\
        );

    \I__7933\ : CascadeMux
    port map (
            O => \N__37640\,
            I => \elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_\
        );

    \I__7932\ : CascadeMux
    port map (
            O => \N__37637\,
            I => \N__37634\
        );

    \I__7931\ : InMux
    port map (
            O => \N__37634\,
            I => \N__37631\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__37631\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__7929\ : IoInMux
    port map (
            O => \N__37628\,
            I => \N__37625\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__37625\,
            I => \N__37622\
        );

    \I__7927\ : IoSpan4Mux
    port map (
            O => \N__37622\,
            I => \N__37619\
        );

    \I__7926\ : Sp12to4
    port map (
            O => \N__37619\,
            I => \N__37616\
        );

    \I__7925\ : Odrv12
    port map (
            O => \N__37616\,
            I => \current_shift_inst.timer_s1.N_166_i\
        );

    \I__7924\ : IoInMux
    port map (
            O => \N__37613\,
            I => \N__37610\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__37610\,
            I => \N__37607\
        );

    \I__7922\ : IoSpan4Mux
    port map (
            O => \N__37607\,
            I => \N__37604\
        );

    \I__7921\ : Span4Mux_s1_v
    port map (
            O => \N__37604\,
            I => \N__37601\
        );

    \I__7920\ : Span4Mux_v
    port map (
            O => \N__37601\,
            I => \N__37596\
        );

    \I__7919\ : InMux
    port map (
            O => \N__37600\,
            I => \N__37591\
        );

    \I__7918\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37591\
        );

    \I__7917\ : Odrv4
    port map (
            O => \N__37596\,
            I => s1_phy_c
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__37591\,
            I => s1_phy_c
        );

    \I__7915\ : InMux
    port map (
            O => \N__37586\,
            I => \N__37582\
        );

    \I__7914\ : InMux
    port map (
            O => \N__37585\,
            I => \N__37579\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__37582\,
            I => \N__37576\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__37579\,
            I => \N__37573\
        );

    \I__7911\ : Span4Mux_h
    port map (
            O => \N__37576\,
            I => \N__37568\
        );

    \I__7910\ : Span4Mux_h
    port map (
            O => \N__37573\,
            I => \N__37568\
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__37568\,
            I => state_ns_i_a3_1
        );

    \I__7908\ : CascadeMux
    port map (
            O => \N__37565\,
            I => \N__37562\
        );

    \I__7907\ : InMux
    port map (
            O => \N__37562\,
            I => \N__37559\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__37559\,
            I => \N__37556\
        );

    \I__7905\ : Span4Mux_v
    port map (
            O => \N__37556\,
            I => \N__37553\
        );

    \I__7904\ : Span4Mux_v
    port map (
            O => \N__37553\,
            I => \N__37548\
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__37552\,
            I => \N__37544\
        );

    \I__7902\ : InMux
    port map (
            O => \N__37551\,
            I => \N__37539\
        );

    \I__7901\ : Span4Mux_h
    port map (
            O => \N__37548\,
            I => \N__37536\
        );

    \I__7900\ : InMux
    port map (
            O => \N__37547\,
            I => \N__37527\
        );

    \I__7899\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37527\
        );

    \I__7898\ : InMux
    port map (
            O => \N__37543\,
            I => \N__37527\
        );

    \I__7897\ : InMux
    port map (
            O => \N__37542\,
            I => \N__37527\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__37539\,
            I => state_3
        );

    \I__7895\ : Odrv4
    port map (
            O => \N__37536\,
            I => state_3
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__37527\,
            I => state_3
        );

    \I__7893\ : InMux
    port map (
            O => \N__37520\,
            I => \N__37515\
        );

    \I__7892\ : InMux
    port map (
            O => \N__37519\,
            I => \N__37512\
        );

    \I__7891\ : InMux
    port map (
            O => \N__37518\,
            I => \N__37509\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__37515\,
            I => \N__37506\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__37512\,
            I => \N__37501\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__37509\,
            I => \N__37501\
        );

    \I__7887\ : Span4Mux_v
    port map (
            O => \N__37506\,
            I => \N__37496\
        );

    \I__7886\ : Span4Mux_v
    port map (
            O => \N__37501\,
            I => \N__37496\
        );

    \I__7885\ : Span4Mux_v
    port map (
            O => \N__37496\,
            I => \N__37493\
        );

    \I__7884\ : Span4Mux_v
    port map (
            O => \N__37493\,
            I => \N__37490\
        );

    \I__7883\ : Span4Mux_v
    port map (
            O => \N__37490\,
            I => \N__37487\
        );

    \I__7882\ : Odrv4
    port map (
            O => \N__37487\,
            I => \il_max_comp1_D2\
        );

    \I__7881\ : InMux
    port map (
            O => \N__37484\,
            I => \N__37481\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__37481\,
            I => \N__37478\
        );

    \I__7879\ : Span4Mux_v
    port map (
            O => \N__37478\,
            I => \N__37475\
        );

    \I__7878\ : Span4Mux_v
    port map (
            O => \N__37475\,
            I => \N__37472\
        );

    \I__7877\ : Odrv4
    port map (
            O => \N__37472\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__7876\ : InMux
    port map (
            O => \N__37469\,
            I => \N__37466\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__37466\,
            I => \N__37463\
        );

    \I__7874\ : Span4Mux_v
    port map (
            O => \N__37463\,
            I => \N__37460\
        );

    \I__7873\ : Span4Mux_v
    port map (
            O => \N__37460\,
            I => \N__37456\
        );

    \I__7872\ : CascadeMux
    port map (
            O => \N__37459\,
            I => \N__37453\
        );

    \I__7871\ : Span4Mux_v
    port map (
            O => \N__37456\,
            I => \N__37448\
        );

    \I__7870\ : InMux
    port map (
            O => \N__37453\,
            I => \N__37443\
        );

    \I__7869\ : InMux
    port map (
            O => \N__37452\,
            I => \N__37443\
        );

    \I__7868\ : InMux
    port map (
            O => \N__37451\,
            I => \N__37440\
        );

    \I__7867\ : Odrv4
    port map (
            O => \N__37448\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__37443\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__37440\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__7864\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37430\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__37430\,
            I => \N__37427\
        );

    \I__7862\ : Span4Mux_v
    port map (
            O => \N__37427\,
            I => \N__37424\
        );

    \I__7861\ : Span4Mux_v
    port map (
            O => \N__37424\,
            I => \N__37420\
        );

    \I__7860\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37415\
        );

    \I__7859\ : Span4Mux_v
    port map (
            O => \N__37420\,
            I => \N__37412\
        );

    \I__7858\ : InMux
    port map (
            O => \N__37419\,
            I => \N__37409\
        );

    \I__7857\ : InMux
    port map (
            O => \N__37418\,
            I => \N__37406\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__37415\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7855\ : Odrv4
    port map (
            O => \N__37412\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__37409\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37406\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7852\ : InMux
    port map (
            O => \N__37397\,
            I => \N__37394\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__37394\,
            I => \N__37389\
        );

    \I__7850\ : CascadeMux
    port map (
            O => \N__37393\,
            I => \N__37386\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37392\,
            I => \N__37383\
        );

    \I__7848\ : Span4Mux_h
    port map (
            O => \N__37389\,
            I => \N__37380\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37386\,
            I => \N__37377\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__37383\,
            I => \N__37374\
        );

    \I__7845\ : Odrv4
    port map (
            O => \N__37380\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__37377\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__7843\ : Odrv4
    port map (
            O => \N__37374\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__7842\ : InMux
    port map (
            O => \N__37367\,
            I => \N__37364\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__37364\,
            I => \N__37361\
        );

    \I__7840\ : Odrv4
    port map (
            O => \N__37361\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37355\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7837\ : Odrv4
    port map (
            O => \N__37352\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__7836\ : InMux
    port map (
            O => \N__37349\,
            I => \N__37346\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__37346\,
            I => \N__37343\
        );

    \I__7834\ : Odrv4
    port map (
            O => \N__37343\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__7833\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37334\
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__37334\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37331\,
            I => \N__37328\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__37328\,
            I => \N__37325\
        );

    \I__7828\ : Odrv4
    port map (
            O => \N__37325\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37319\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__37319\,
            I => \N__37316\
        );

    \I__7825\ : Odrv12
    port map (
            O => \N__37316\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__7824\ : CascadeMux
    port map (
            O => \N__37313\,
            I => \N__37310\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37310\,
            I => \N__37307\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__37307\,
            I => \N__37304\
        );

    \I__7821\ : Odrv4
    port map (
            O => \N__37304\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__7820\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37298\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__37298\,
            I => \N__37295\
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__37295\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__7817\ : InMux
    port map (
            O => \N__37292\,
            I => \N__37289\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__37289\,
            I => \N__37286\
        );

    \I__7815\ : Odrv12
    port map (
            O => \N__37286\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37280\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__37280\,
            I => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37274\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__37274\,
            I => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\
        );

    \I__7810\ : CascadeMux
    port map (
            O => \N__37271\,
            I => \N__37268\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37268\,
            I => \N__37265\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__37265\,
            I => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37259\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__37259\,
            I => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\
        );

    \I__7805\ : CascadeMux
    port map (
            O => \N__37256\,
            I => \N__37253\
        );

    \I__7804\ : InMux
    port map (
            O => \N__37253\,
            I => \N__37247\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37247\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__37247\,
            I => \N__37244\
        );

    \I__7801\ : Span4Mux_h
    port map (
            O => \N__37244\,
            I => \N__37240\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37243\,
            I => \N__37237\
        );

    \I__7799\ : Span4Mux_h
    port map (
            O => \N__37240\,
            I => \N__37234\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__37237\,
            I => \elapsed_time_ns_1_RNI81DJ11_0_2\
        );

    \I__7797\ : Odrv4
    port map (
            O => \N__37234\,
            I => \elapsed_time_ns_1_RNI81DJ11_0_2\
        );

    \I__7796\ : InMux
    port map (
            O => \N__37229\,
            I => \N__37226\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__37226\,
            I => \N__37222\
        );

    \I__7794\ : InMux
    port map (
            O => \N__37225\,
            I => \N__37219\
        );

    \I__7793\ : Span4Mux_v
    port map (
            O => \N__37222\,
            I => \N__37215\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37219\,
            I => \N__37212\
        );

    \I__7791\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37209\
        );

    \I__7790\ : Odrv4
    port map (
            O => \N__37215\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__7789\ : Odrv12
    port map (
            O => \N__37212\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__37209\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37195\
        );

    \I__7786\ : InMux
    port map (
            O => \N__37201\,
            I => \N__37195\
        );

    \I__7785\ : CascadeMux
    port map (
            O => \N__37200\,
            I => \N__37192\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__37195\,
            I => \N__37189\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37192\,
            I => \N__37186\
        );

    \I__7782\ : Span4Mux_h
    port map (
            O => \N__37189\,
            I => \N__37183\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__37186\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__7780\ : Odrv4
    port map (
            O => \N__37183\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__7779\ : CEMux
    port map (
            O => \N__37178\,
            I => \N__37163\
        );

    \I__7778\ : CEMux
    port map (
            O => \N__37177\,
            I => \N__37163\
        );

    \I__7777\ : CEMux
    port map (
            O => \N__37176\,
            I => \N__37163\
        );

    \I__7776\ : CEMux
    port map (
            O => \N__37175\,
            I => \N__37163\
        );

    \I__7775\ : CEMux
    port map (
            O => \N__37174\,
            I => \N__37163\
        );

    \I__7774\ : GlobalMux
    port map (
            O => \N__37163\,
            I => \N__37160\
        );

    \I__7773\ : gio2CtrlBuf
    port map (
            O => \N__37160\,
            I => \delay_measurement_inst.delay_hc_timer.N_432_i_g\
        );

    \I__7772\ : InMux
    port map (
            O => \N__37157\,
            I => \N__37148\
        );

    \I__7771\ : InMux
    port map (
            O => \N__37156\,
            I => \N__37148\
        );

    \I__7770\ : CascadeMux
    port map (
            O => \N__37155\,
            I => \N__37138\
        );

    \I__7769\ : InMux
    port map (
            O => \N__37154\,
            I => \N__37135\
        );

    \I__7768\ : CascadeMux
    port map (
            O => \N__37153\,
            I => \N__37132\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__37148\,
            I => \N__37128\
        );

    \I__7766\ : InMux
    port map (
            O => \N__37147\,
            I => \N__37125\
        );

    \I__7765\ : InMux
    port map (
            O => \N__37146\,
            I => \N__37122\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37145\,
            I => \N__37119\
        );

    \I__7763\ : InMux
    port map (
            O => \N__37144\,
            I => \N__37116\
        );

    \I__7762\ : InMux
    port map (
            O => \N__37143\,
            I => \N__37107\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37142\,
            I => \N__37107\
        );

    \I__7760\ : InMux
    port map (
            O => \N__37141\,
            I => \N__37107\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37138\,
            I => \N__37107\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__37135\,
            I => \N__37099\
        );

    \I__7757\ : InMux
    port map (
            O => \N__37132\,
            I => \N__37096\
        );

    \I__7756\ : InMux
    port map (
            O => \N__37131\,
            I => \N__37093\
        );

    \I__7755\ : Span4Mux_h
    port map (
            O => \N__37128\,
            I => \N__37090\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__37125\,
            I => \N__37079\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__37122\,
            I => \N__37079\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__37119\,
            I => \N__37079\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__37116\,
            I => \N__37079\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__37107\,
            I => \N__37079\
        );

    \I__7749\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37072\
        );

    \I__7748\ : InMux
    port map (
            O => \N__37105\,
            I => \N__37069\
        );

    \I__7747\ : InMux
    port map (
            O => \N__37104\,
            I => \N__37066\
        );

    \I__7746\ : InMux
    port map (
            O => \N__37103\,
            I => \N__37061\
        );

    \I__7745\ : InMux
    port map (
            O => \N__37102\,
            I => \N__37061\
        );

    \I__7744\ : Span4Mux_h
    port map (
            O => \N__37099\,
            I => \N__37058\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__37096\,
            I => \N__37049\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__37093\,
            I => \N__37049\
        );

    \I__7741\ : Span4Mux_v
    port map (
            O => \N__37090\,
            I => \N__37049\
        );

    \I__7740\ : Span4Mux_v
    port map (
            O => \N__37079\,
            I => \N__37049\
        );

    \I__7739\ : InMux
    port map (
            O => \N__37078\,
            I => \N__37040\
        );

    \I__7738\ : InMux
    port map (
            O => \N__37077\,
            I => \N__37040\
        );

    \I__7737\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37040\
        );

    \I__7736\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37040\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__37072\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__37069\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__37066\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__37061\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__37058\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__37049\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__37040\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\
        );

    \I__7728\ : CascadeMux
    port map (
            O => \N__37025\,
            I => \N__37022\
        );

    \I__7727\ : InMux
    port map (
            O => \N__37022\,
            I => \N__37019\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__37019\,
            I => \N__37015\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__37018\,
            I => \N__37012\
        );

    \I__7724\ : Span12Mux_h
    port map (
            O => \N__37015\,
            I => \N__37009\
        );

    \I__7723\ : InMux
    port map (
            O => \N__37012\,
            I => \N__37006\
        );

    \I__7722\ : Odrv12
    port map (
            O => \N__37009\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__37006\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__7720\ : InMux
    port map (
            O => \N__37001\,
            I => \N__36991\
        );

    \I__7719\ : CascadeMux
    port map (
            O => \N__37000\,
            I => \N__36988\
        );

    \I__7718\ : CascadeMux
    port map (
            O => \N__36999\,
            I => \N__36985\
        );

    \I__7717\ : InMux
    port map (
            O => \N__36998\,
            I => \N__36975\
        );

    \I__7716\ : InMux
    port map (
            O => \N__36997\,
            I => \N__36975\
        );

    \I__7715\ : CascadeMux
    port map (
            O => \N__36996\,
            I => \N__36971\
        );

    \I__7714\ : CascadeMux
    port map (
            O => \N__36995\,
            I => \N__36966\
        );

    \I__7713\ : CascadeMux
    port map (
            O => \N__36994\,
            I => \N__36963\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__36991\,
            I => \N__36958\
        );

    \I__7711\ : InMux
    port map (
            O => \N__36988\,
            I => \N__36953\
        );

    \I__7710\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36953\
        );

    \I__7709\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36948\
        );

    \I__7708\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36948\
        );

    \I__7707\ : CascadeMux
    port map (
            O => \N__36982\,
            I => \N__36945\
        );

    \I__7706\ : InMux
    port map (
            O => \N__36981\,
            I => \N__36941\
        );

    \I__7705\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36938\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__36975\,
            I => \N__36935\
        );

    \I__7703\ : InMux
    port map (
            O => \N__36974\,
            I => \N__36929\
        );

    \I__7702\ : InMux
    port map (
            O => \N__36971\,
            I => \N__36929\
        );

    \I__7701\ : InMux
    port map (
            O => \N__36970\,
            I => \N__36926\
        );

    \I__7700\ : InMux
    port map (
            O => \N__36969\,
            I => \N__36921\
        );

    \I__7699\ : InMux
    port map (
            O => \N__36966\,
            I => \N__36921\
        );

    \I__7698\ : InMux
    port map (
            O => \N__36963\,
            I => \N__36918\
        );

    \I__7697\ : InMux
    port map (
            O => \N__36962\,
            I => \N__36913\
        );

    \I__7696\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36913\
        );

    \I__7695\ : Span4Mux_h
    port map (
            O => \N__36958\,
            I => \N__36906\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__36953\,
            I => \N__36906\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__36948\,
            I => \N__36906\
        );

    \I__7692\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36903\
        );

    \I__7691\ : InMux
    port map (
            O => \N__36944\,
            I => \N__36900\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__36941\,
            I => \N__36892\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__36938\,
            I => \N__36887\
        );

    \I__7688\ : Span4Mux_h
    port map (
            O => \N__36935\,
            I => \N__36887\
        );

    \I__7687\ : InMux
    port map (
            O => \N__36934\,
            I => \N__36884\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__36929\,
            I => \N__36869\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__36926\,
            I => \N__36869\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__36921\,
            I => \N__36869\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__36918\,
            I => \N__36869\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__36913\,
            I => \N__36869\
        );

    \I__7681\ : Span4Mux_h
    port map (
            O => \N__36906\,
            I => \N__36869\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__36903\,
            I => \N__36869\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__36900\,
            I => \N__36861\
        );

    \I__7678\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36856\
        );

    \I__7677\ : InMux
    port map (
            O => \N__36898\,
            I => \N__36856\
        );

    \I__7676\ : InMux
    port map (
            O => \N__36897\,
            I => \N__36849\
        );

    \I__7675\ : InMux
    port map (
            O => \N__36896\,
            I => \N__36849\
        );

    \I__7674\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36849\
        );

    \I__7673\ : Span4Mux_v
    port map (
            O => \N__36892\,
            I => \N__36840\
        );

    \I__7672\ : Span4Mux_v
    port map (
            O => \N__36887\,
            I => \N__36840\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__36884\,
            I => \N__36840\
        );

    \I__7670\ : Span4Mux_v
    port map (
            O => \N__36869\,
            I => \N__36840\
        );

    \I__7669\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36829\
        );

    \I__7668\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36829\
        );

    \I__7667\ : InMux
    port map (
            O => \N__36866\,
            I => \N__36829\
        );

    \I__7666\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36829\
        );

    \I__7665\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36829\
        );

    \I__7664\ : Span4Mux_h
    port map (
            O => \N__36861\,
            I => \N__36826\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__36856\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__36849\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__36840\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__36829\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__7659\ : Odrv4
    port map (
            O => \N__36826\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i\
        );

    \I__7658\ : InMux
    port map (
            O => \N__36815\,
            I => \N__36812\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__36812\,
            I => \N__36809\
        );

    \I__7656\ : Span4Mux_h
    port map (
            O => \N__36809\,
            I => \N__36805\
        );

    \I__7655\ : InMux
    port map (
            O => \N__36808\,
            I => \N__36802\
        );

    \I__7654\ : Span4Mux_h
    port map (
            O => \N__36805\,
            I => \N__36799\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__36802\,
            I => \elapsed_time_ns_1_RNIO1ND11_0_20\
        );

    \I__7652\ : Odrv4
    port map (
            O => \N__36799\,
            I => \elapsed_time_ns_1_RNIO1ND11_0_20\
        );

    \I__7651\ : InMux
    port map (
            O => \N__36794\,
            I => \N__36791\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__36791\,
            I => \N__36788\
        );

    \I__7649\ : Odrv4
    port map (
            O => \N__36788\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__7648\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36782\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__36782\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__7646\ : InMux
    port map (
            O => \N__36779\,
            I => \N__36776\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__36776\,
            I => \N__36773\
        );

    \I__7644\ : Span4Mux_h
    port map (
            O => \N__36773\,
            I => \N__36770\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__36770\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__7642\ : InMux
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__36764\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__7640\ : InMux
    port map (
            O => \N__36761\,
            I => \N__36758\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__36758\,
            I => \N__36755\
        );

    \I__7638\ : Odrv4
    port map (
            O => \N__36755\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__7637\ : InMux
    port map (
            O => \N__36752\,
            I => \N__36749\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__36749\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__36746\,
            I => \N__36743\
        );

    \I__7634\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36740\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__36740\,
            I => \N__36737\
        );

    \I__7632\ : Odrv4
    port map (
            O => \N__36737\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__7631\ : InMux
    port map (
            O => \N__36734\,
            I => \N__36731\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__36731\,
            I => \N__36728\
        );

    \I__7629\ : Odrv4
    port map (
            O => \N__36728\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__7628\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36722\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__36722\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__7626\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36716\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__36716\,
            I => \N__36713\
        );

    \I__7624\ : Span4Mux_h
    port map (
            O => \N__36713\,
            I => \N__36710\
        );

    \I__7623\ : Odrv4
    port map (
            O => \N__36710\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__7622\ : InMux
    port map (
            O => \N__36707\,
            I => \N__36704\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__36704\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__7620\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36698\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__36698\,
            I => \N__36695\
        );

    \I__7618\ : Odrv4
    port map (
            O => \N__36695\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__7617\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36689\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36686\
        );

    \I__7615\ : Odrv12
    port map (
            O => \N__36686\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__7614\ : InMux
    port map (
            O => \N__36683\,
            I => \N__36680\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__36680\,
            I => \N__36677\
        );

    \I__7612\ : Odrv4
    port map (
            O => \N__36677\,
            I => \current_shift_inst.control_input_1_axb_11\
        );

    \I__7611\ : InMux
    port map (
            O => \N__36674\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__7610\ : InMux
    port map (
            O => \N__36671\,
            I => \N__36668\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__36668\,
            I => \N__36665\
        );

    \I__7608\ : Span4Mux_v
    port map (
            O => \N__36665\,
            I => \N__36661\
        );

    \I__7607\ : InMux
    port map (
            O => \N__36664\,
            I => \N__36658\
        );

    \I__7606\ : Span4Mux_v
    port map (
            O => \N__36661\,
            I => \N__36653\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__36658\,
            I => \N__36653\
        );

    \I__7604\ : Odrv4
    port map (
            O => \N__36653\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__7603\ : CascadeMux
    port map (
            O => \N__36650\,
            I => \N__36647\
        );

    \I__7602\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36644\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__36644\,
            I => \N__36641\
        );

    \I__7600\ : Odrv4
    port map (
            O => \N__36641\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__7599\ : CascadeMux
    port map (
            O => \N__36638\,
            I => \N__36634\
        );

    \I__7598\ : InMux
    port map (
            O => \N__36637\,
            I => \N__36631\
        );

    \I__7597\ : InMux
    port map (
            O => \N__36634\,
            I => \N__36628\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__36631\,
            I => \current_shift_inst.N_1609_i\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__36628\,
            I => \current_shift_inst.N_1609_i\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__36623\,
            I => \N__36620\
        );

    \I__7593\ : InMux
    port map (
            O => \N__36620\,
            I => \N__36617\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__36617\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__7591\ : InMux
    port map (
            O => \N__36614\,
            I => \N__36611\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__36611\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__7589\ : InMux
    port map (
            O => \N__36608\,
            I => \N__36605\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__36605\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__7587\ : InMux
    port map (
            O => \N__36602\,
            I => \N__36599\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__36599\,
            I => \N__36596\
        );

    \I__7585\ : Odrv4
    port map (
            O => \N__36596\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__7584\ : InMux
    port map (
            O => \N__36593\,
            I => \N__36590\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__36590\,
            I => \N__36587\
        );

    \I__7582\ : Odrv4
    port map (
            O => \N__36587\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__7581\ : InMux
    port map (
            O => \N__36584\,
            I => \N__36581\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__36581\,
            I => \N__36578\
        );

    \I__7579\ : Span4Mux_v
    port map (
            O => \N__36578\,
            I => \N__36575\
        );

    \I__7578\ : Odrv4
    port map (
            O => \N__36575\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__7577\ : InMux
    port map (
            O => \N__36572\,
            I => \N__36569\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__36569\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__7575\ : InMux
    port map (
            O => \N__36566\,
            I => \N__36563\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__36563\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__7573\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36557\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__36557\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__7571\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36551\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__36551\,
            I => \N__36548\
        );

    \I__7569\ : Span4Mux_v
    port map (
            O => \N__36548\,
            I => \N__36545\
        );

    \I__7568\ : Odrv4
    port map (
            O => \N__36545\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__7567\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36539\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__36539\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__7565\ : InMux
    port map (
            O => \N__36536\,
            I => \N__36533\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__36533\,
            I => \N__36530\
        );

    \I__7563\ : Span4Mux_h
    port map (
            O => \N__36530\,
            I => \N__36527\
        );

    \I__7562\ : Odrv4
    port map (
            O => \N__36527\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__7561\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36521\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__36521\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__7559\ : InMux
    port map (
            O => \N__36518\,
            I => \N__36515\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__36515\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__7557\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36509\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__36509\,
            I => \N__36506\
        );

    \I__7555\ : Span4Mux_v
    port map (
            O => \N__36506\,
            I => \N__36503\
        );

    \I__7554\ : Odrv4
    port map (
            O => \N__36503\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__7553\ : InMux
    port map (
            O => \N__36500\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__7552\ : InMux
    port map (
            O => \N__36497\,
            I => \N__36494\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__36494\,
            I => \N__36491\
        );

    \I__7550\ : Span4Mux_h
    port map (
            O => \N__36491\,
            I => \N__36488\
        );

    \I__7549\ : Odrv4
    port map (
            O => \N__36488\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__7548\ : InMux
    port map (
            O => \N__36485\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__7547\ : InMux
    port map (
            O => \N__36482\,
            I => \N__36479\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36476\
        );

    \I__7545\ : Span4Mux_v
    port map (
            O => \N__36476\,
            I => \N__36473\
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__36473\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__7543\ : InMux
    port map (
            O => \N__36470\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__7542\ : InMux
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__36464\,
            I => \N__36461\
        );

    \I__7540\ : Span4Mux_h
    port map (
            O => \N__36461\,
            I => \N__36458\
        );

    \I__7539\ : Odrv4
    port map (
            O => \N__36458\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__7538\ : InMux
    port map (
            O => \N__36455\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36452\,
            I => \N__36449\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__36449\,
            I => \N__36446\
        );

    \I__7535\ : Span4Mux_v
    port map (
            O => \N__36446\,
            I => \N__36443\
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__36443\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__7533\ : InMux
    port map (
            O => \N__36440\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__7532\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36434\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__36434\,
            I => \N__36431\
        );

    \I__7530\ : Span4Mux_h
    port map (
            O => \N__36431\,
            I => \N__36428\
        );

    \I__7529\ : Odrv4
    port map (
            O => \N__36428\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36425\,
            I => \bfn_15_17_0_\
        );

    \I__7527\ : InMux
    port map (
            O => \N__36422\,
            I => \N__36419\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__36419\,
            I => \N__36416\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__36416\,
            I => \N__36413\
        );

    \I__7524\ : Odrv4
    port map (
            O => \N__36413\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__7523\ : InMux
    port map (
            O => \N__36410\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__7522\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36404\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__36404\,
            I => \N__36401\
        );

    \I__7520\ : Span4Mux_v
    port map (
            O => \N__36401\,
            I => \N__36398\
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__36398\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36395\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36392\,
            I => \N__36388\
        );

    \I__7516\ : InMux
    port map (
            O => \N__36391\,
            I => \N__36385\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__36388\,
            I => \N__36382\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__36385\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__7513\ : Odrv12
    port map (
            O => \N__36382\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__7512\ : InMux
    port map (
            O => \N__36377\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__7511\ : InMux
    port map (
            O => \N__36374\,
            I => \N__36370\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36373\,
            I => \N__36367\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__36370\,
            I => \N__36364\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__36367\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7507\ : Odrv4
    port map (
            O => \N__36364\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7506\ : InMux
    port map (
            O => \N__36359\,
            I => \bfn_15_15_0_\
        );

    \I__7505\ : InMux
    port map (
            O => \N__36356\,
            I => \N__36352\
        );

    \I__7504\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36349\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__36352\,
            I => \N__36346\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__36349\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7501\ : Odrv4
    port map (
            O => \N__36346\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36341\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36338\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__7498\ : InMux
    port map (
            O => \N__36335\,
            I => \N__36331\
        );

    \I__7497\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36328\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__36331\,
            I => \N__36325\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__36328\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7494\ : Odrv4
    port map (
            O => \N__36325\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7493\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36317\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__36317\,
            I => \N__36314\
        );

    \I__7491\ : Span12Mux_v
    port map (
            O => \N__36314\,
            I => \N__36311\
        );

    \I__7490\ : Odrv12
    port map (
            O => \N__36311\,
            I => \phase_controller_inst1.stoper_hc.un1_start_latched2_0\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36308\,
            I => \N__36305\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__36305\,
            I => \N__36302\
        );

    \I__7487\ : Span4Mux_v
    port map (
            O => \N__36302\,
            I => \N__36297\
        );

    \I__7486\ : InMux
    port map (
            O => \N__36301\,
            I => \N__36294\
        );

    \I__7485\ : CascadeMux
    port map (
            O => \N__36300\,
            I => \N__36290\
        );

    \I__7484\ : Span4Mux_h
    port map (
            O => \N__36297\,
            I => \N__36285\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__36294\,
            I => \N__36285\
        );

    \I__7482\ : CascadeMux
    port map (
            O => \N__36293\,
            I => \N__36281\
        );

    \I__7481\ : InMux
    port map (
            O => \N__36290\,
            I => \N__36276\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__36285\,
            I => \N__36273\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36284\,
            I => \N__36270\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36281\,
            I => \N__36263\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36280\,
            I => \N__36263\
        );

    \I__7476\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36263\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__36276\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__36273\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__36270\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__36263\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7471\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36248\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36245\
        );

    \I__7469\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36242\
        );

    \I__7468\ : CascadeMux
    port map (
            O => \N__36251\,
            I => \N__36236\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__36248\,
            I => \N__36233\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__36245\,
            I => \N__36228\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__36242\,
            I => \N__36228\
        );

    \I__7464\ : InMux
    port map (
            O => \N__36241\,
            I => \N__36221\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36240\,
            I => \N__36221\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36239\,
            I => \N__36221\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36217\
        );

    \I__7460\ : Span4Mux_v
    port map (
            O => \N__36233\,
            I => \N__36214\
        );

    \I__7459\ : Sp12to4
    port map (
            O => \N__36228\,
            I => \N__36209\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36221\,
            I => \N__36209\
        );

    \I__7457\ : InMux
    port map (
            O => \N__36220\,
            I => \N__36206\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__36217\,
            I => \N__36203\
        );

    \I__7455\ : Sp12to4
    port map (
            O => \N__36214\,
            I => \N__36198\
        );

    \I__7454\ : Span12Mux_v
    port map (
            O => \N__36209\,
            I => \N__36198\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__36206\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7452\ : Odrv4
    port map (
            O => \N__36203\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7451\ : Odrv12
    port map (
            O => \N__36198\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36186\
        );

    \I__7449\ : InMux
    port map (
            O => \N__36190\,
            I => \N__36181\
        );

    \I__7448\ : InMux
    port map (
            O => \N__36189\,
            I => \N__36181\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__36186\,
            I => \N__36177\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__36181\,
            I => \N__36174\
        );

    \I__7445\ : InMux
    port map (
            O => \N__36180\,
            I => \N__36171\
        );

    \I__7444\ : Span4Mux_v
    port map (
            O => \N__36177\,
            I => \N__36166\
        );

    \I__7443\ : Span4Mux_h
    port map (
            O => \N__36174\,
            I => \N__36166\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__36171\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__7441\ : Odrv4
    port map (
            O => \N__36166\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__7440\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36158\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__36158\,
            I => \N__36154\
        );

    \I__7438\ : InMux
    port map (
            O => \N__36157\,
            I => \N__36151\
        );

    \I__7437\ : Span4Mux_v
    port map (
            O => \N__36154\,
            I => \N__36146\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36151\,
            I => \N__36146\
        );

    \I__7435\ : Span4Mux_v
    port map (
            O => \N__36146\,
            I => \N__36143\
        );

    \I__7434\ : Span4Mux_h
    port map (
            O => \N__36143\,
            I => \N__36140\
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__36140\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__7432\ : InMux
    port map (
            O => \N__36137\,
            I => \N__36134\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__36134\,
            I => \N__36131\
        );

    \I__7430\ : Odrv12
    port map (
            O => \N__36131\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36128\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36122\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__36122\,
            I => \N__36119\
        );

    \I__7426\ : Span4Mux_h
    port map (
            O => \N__36119\,
            I => \N__36116\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__36116\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36113\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__7423\ : InMux
    port map (
            O => \N__36110\,
            I => \N__36106\
        );

    \I__7422\ : InMux
    port map (
            O => \N__36109\,
            I => \N__36103\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__36106\,
            I => \N__36100\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__36103\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7419\ : Odrv12
    port map (
            O => \N__36100\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7418\ : InMux
    port map (
            O => \N__36095\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__7417\ : InMux
    port map (
            O => \N__36092\,
            I => \N__36088\
        );

    \I__7416\ : InMux
    port map (
            O => \N__36091\,
            I => \N__36085\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__36088\,
            I => \N__36082\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__36085\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7413\ : Odrv12
    port map (
            O => \N__36082\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7412\ : InMux
    port map (
            O => \N__36077\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36074\,
            I => \N__36070\
        );

    \I__7410\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36067\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__36070\,
            I => \N__36064\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__36067\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7407\ : Odrv4
    port map (
            O => \N__36064\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7406\ : InMux
    port map (
            O => \N__36059\,
            I => \bfn_15_14_0_\
        );

    \I__7405\ : InMux
    port map (
            O => \N__36056\,
            I => \N__36052\
        );

    \I__7404\ : InMux
    port map (
            O => \N__36055\,
            I => \N__36049\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__36052\,
            I => \N__36046\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__36049\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7401\ : Odrv4
    port map (
            O => \N__36046\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7400\ : InMux
    port map (
            O => \N__36041\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36038\,
            I => \N__36034\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36031\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__36034\,
            I => \N__36028\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__36031\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7395\ : Odrv4
    port map (
            O => \N__36028\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7394\ : InMux
    port map (
            O => \N__36023\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__7393\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36016\
        );

    \I__7392\ : InMux
    port map (
            O => \N__36019\,
            I => \N__36013\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__36016\,
            I => \N__36010\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__36013\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__36010\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7388\ : InMux
    port map (
            O => \N__36005\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__7387\ : InMux
    port map (
            O => \N__36002\,
            I => \N__35999\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__35999\,
            I => \N__35995\
        );

    \I__7385\ : InMux
    port map (
            O => \N__35998\,
            I => \N__35992\
        );

    \I__7384\ : Span4Mux_v
    port map (
            O => \N__35995\,
            I => \N__35989\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__35992\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7382\ : Odrv4
    port map (
            O => \N__35989\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7381\ : InMux
    port map (
            O => \N__35984\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__7380\ : InMux
    port map (
            O => \N__35981\,
            I => \N__35977\
        );

    \I__7379\ : InMux
    port map (
            O => \N__35980\,
            I => \N__35974\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__35977\,
            I => \N__35971\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__35974\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7376\ : Odrv4
    port map (
            O => \N__35971\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7375\ : InMux
    port map (
            O => \N__35966\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__7374\ : InMux
    port map (
            O => \N__35963\,
            I => \N__35960\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__35960\,
            I => \N__35956\
        );

    \I__7372\ : InMux
    port map (
            O => \N__35959\,
            I => \N__35953\
        );

    \I__7371\ : Span4Mux_v
    port map (
            O => \N__35956\,
            I => \N__35950\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__35953\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7369\ : Odrv4
    port map (
            O => \N__35950\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7368\ : InMux
    port map (
            O => \N__35945\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__7367\ : InMux
    port map (
            O => \N__35942\,
            I => \N__35939\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__35939\,
            I => \N__35936\
        );

    \I__7365\ : Span4Mux_h
    port map (
            O => \N__35936\,
            I => \N__35933\
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__35933\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__7363\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35923\
        );

    \I__7362\ : InMux
    port map (
            O => \N__35929\,
            I => \N__35919\
        );

    \I__7361\ : InMux
    port map (
            O => \N__35928\,
            I => \N__35914\
        );

    \I__7360\ : InMux
    port map (
            O => \N__35927\,
            I => \N__35911\
        );

    \I__7359\ : InMux
    port map (
            O => \N__35926\,
            I => \N__35908\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__35923\,
            I => \N__35905\
        );

    \I__7357\ : CascadeMux
    port map (
            O => \N__35922\,
            I => \N__35902\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__35919\,
            I => \N__35899\
        );

    \I__7355\ : InMux
    port map (
            O => \N__35918\,
            I => \N__35894\
        );

    \I__7354\ : InMux
    port map (
            O => \N__35917\,
            I => \N__35894\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__35914\,
            I => \N__35891\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__35911\,
            I => \N__35886\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__35908\,
            I => \N__35886\
        );

    \I__7350\ : Span4Mux_v
    port map (
            O => \N__35905\,
            I => \N__35883\
        );

    \I__7349\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35880\
        );

    \I__7348\ : Span4Mux_v
    port map (
            O => \N__35899\,
            I => \N__35877\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__35894\,
            I => \N__35874\
        );

    \I__7346\ : Span4Mux_v
    port map (
            O => \N__35891\,
            I => \N__35867\
        );

    \I__7345\ : Span4Mux_v
    port map (
            O => \N__35886\,
            I => \N__35867\
        );

    \I__7344\ : Span4Mux_h
    port map (
            O => \N__35883\,
            I => \N__35867\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__35880\,
            I => \N__35862\
        );

    \I__7342\ : Span4Mux_h
    port map (
            O => \N__35877\,
            I => \N__35862\
        );

    \I__7341\ : Odrv12
    port map (
            O => \N__35874\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__35867\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__35862\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5\
        );

    \I__7338\ : CascadeMux
    port map (
            O => \N__35855\,
            I => \N__35852\
        );

    \I__7337\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35849\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__35849\,
            I => \N__35846\
        );

    \I__7335\ : Span4Mux_h
    port map (
            O => \N__35846\,
            I => \N__35840\
        );

    \I__7334\ : InMux
    port map (
            O => \N__35845\,
            I => \N__35837\
        );

    \I__7333\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35834\
        );

    \I__7332\ : InMux
    port map (
            O => \N__35843\,
            I => \N__35831\
        );

    \I__7331\ : Odrv4
    port map (
            O => \N__35840\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__35837\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__35834\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__35831\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\
        );

    \I__7327\ : InMux
    port map (
            O => \N__35822\,
            I => \N__35817\
        );

    \I__7326\ : InMux
    port map (
            O => \N__35821\,
            I => \N__35810\
        );

    \I__7325\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35810\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__35817\,
            I => \N__35807\
        );

    \I__7323\ : CascadeMux
    port map (
            O => \N__35816\,
            I => \N__35804\
        );

    \I__7322\ : InMux
    port map (
            O => \N__35815\,
            I => \N__35801\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__35810\,
            I => \N__35798\
        );

    \I__7320\ : Span4Mux_h
    port map (
            O => \N__35807\,
            I => \N__35795\
        );

    \I__7319\ : InMux
    port map (
            O => \N__35804\,
            I => \N__35792\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__35801\,
            I => \N__35785\
        );

    \I__7317\ : Span4Mux_v
    port map (
            O => \N__35798\,
            I => \N__35785\
        );

    \I__7316\ : Span4Mux_h
    port map (
            O => \N__35795\,
            I => \N__35785\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__35792\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9\
        );

    \I__7314\ : Odrv4
    port map (
            O => \N__35785\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9\
        );

    \I__7313\ : InMux
    port map (
            O => \N__35780\,
            I => \N__35777\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__35777\,
            I => \N__35774\
        );

    \I__7311\ : Span4Mux_v
    port map (
            O => \N__35774\,
            I => \N__35771\
        );

    \I__7310\ : Span4Mux_h
    port map (
            O => \N__35771\,
            I => \N__35768\
        );

    \I__7309\ : Odrv4
    port map (
            O => \N__35768\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\
        );

    \I__7308\ : InMux
    port map (
            O => \N__35765\,
            I => \N__35762\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__35762\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__7306\ : CascadeMux
    port map (
            O => \N__35759\,
            I => \N__35756\
        );

    \I__7305\ : InMux
    port map (
            O => \N__35756\,
            I => \N__35752\
        );

    \I__7304\ : InMux
    port map (
            O => \N__35755\,
            I => \N__35749\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__35752\,
            I => \N__35746\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__35749\,
            I => \N__35743\
        );

    \I__7301\ : Span4Mux_v
    port map (
            O => \N__35746\,
            I => \N__35739\
        );

    \I__7300\ : Span4Mux_h
    port map (
            O => \N__35743\,
            I => \N__35736\
        );

    \I__7299\ : CascadeMux
    port map (
            O => \N__35742\,
            I => \N__35733\
        );

    \I__7298\ : Span4Mux_h
    port map (
            O => \N__35739\,
            I => \N__35728\
        );

    \I__7297\ : Span4Mux_v
    port map (
            O => \N__35736\,
            I => \N__35728\
        );

    \I__7296\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35725\
        );

    \I__7295\ : Span4Mux_h
    port map (
            O => \N__35728\,
            I => \N__35722\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__35725\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7293\ : Odrv4
    port map (
            O => \N__35722\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7292\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35713\
        );

    \I__7291\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35710\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__35713\,
            I => \N__35707\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__35710\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7288\ : Odrv4
    port map (
            O => \N__35707\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7287\ : InMux
    port map (
            O => \N__35702\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__7286\ : CascadeMux
    port map (
            O => \N__35699\,
            I => \N__35696\
        );

    \I__7285\ : InMux
    port map (
            O => \N__35696\,
            I => \N__35693\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__35693\,
            I => \N__35690\
        );

    \I__7283\ : Odrv4
    port map (
            O => \N__35690\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQZ0Z1\
        );

    \I__7282\ : InMux
    port map (
            O => \N__35687\,
            I => \N__35683\
        );

    \I__7281\ : InMux
    port map (
            O => \N__35686\,
            I => \N__35680\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__35683\,
            I => \N__35677\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__35680\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7278\ : Odrv4
    port map (
            O => \N__35677\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7277\ : InMux
    port map (
            O => \N__35672\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__7276\ : InMux
    port map (
            O => \N__35669\,
            I => \N__35665\
        );

    \I__7275\ : InMux
    port map (
            O => \N__35668\,
            I => \N__35662\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__35665\,
            I => \N__35659\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__35662\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7272\ : Odrv4
    port map (
            O => \N__35659\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7271\ : InMux
    port map (
            O => \N__35654\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__7270\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35647\
        );

    \I__7269\ : InMux
    port map (
            O => \N__35650\,
            I => \N__35644\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__35647\,
            I => \N__35641\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__35644\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7266\ : Odrv4
    port map (
            O => \N__35641\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7265\ : InMux
    port map (
            O => \N__35636\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__7264\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35629\
        );

    \I__7263\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35626\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__35629\,
            I => \N__35623\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__35626\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7260\ : Odrv4
    port map (
            O => \N__35623\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7259\ : InMux
    port map (
            O => \N__35618\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__7258\ : CascadeMux
    port map (
            O => \N__35615\,
            I => \N__35612\
        );

    \I__7257\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35609\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__35609\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__7255\ : CascadeMux
    port map (
            O => \N__35606\,
            I => \N__35603\
        );

    \I__7254\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35600\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__35600\,
            I => \N__35597\
        );

    \I__7252\ : Odrv4
    port map (
            O => \N__35597\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__7251\ : CascadeMux
    port map (
            O => \N__35594\,
            I => \N__35591\
        );

    \I__7250\ : InMux
    port map (
            O => \N__35591\,
            I => \N__35588\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__35588\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__7248\ : CascadeMux
    port map (
            O => \N__35585\,
            I => \N__35582\
        );

    \I__7247\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35579\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__35579\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\
        );

    \I__7245\ : CascadeMux
    port map (
            O => \N__35576\,
            I => \N__35573\
        );

    \I__7244\ : InMux
    port map (
            O => \N__35573\,
            I => \N__35570\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__35570\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\
        );

    \I__7242\ : CascadeMux
    port map (
            O => \N__35567\,
            I => \N__35564\
        );

    \I__7241\ : InMux
    port map (
            O => \N__35564\,
            I => \N__35561\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__35561\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\
        );

    \I__7239\ : CascadeMux
    port map (
            O => \N__35558\,
            I => \N__35555\
        );

    \I__7238\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35552\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__35552\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\
        );

    \I__7236\ : InMux
    port map (
            O => \N__35549\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_19\
        );

    \I__7235\ : InMux
    port map (
            O => \N__35546\,
            I => \N__35543\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__35543\,
            I => \N__35540\
        );

    \I__7233\ : Span4Mux_h
    port map (
            O => \N__35540\,
            I => \N__35536\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35533\
        );

    \I__7231\ : Odrv4
    port map (
            O => \N__35536\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__35533\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO\
        );

    \I__7229\ : InMux
    port map (
            O => \N__35528\,
            I => \N__35525\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__35525\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__35522\,
            I => \N__35519\
        );

    \I__7226\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35516\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__35516\,
            I => \N__35513\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__35513\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__7223\ : CascadeMux
    port map (
            O => \N__35510\,
            I => \N__35507\
        );

    \I__7222\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35504\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__35504\,
            I => \N__35501\
        );

    \I__7220\ : Odrv4
    port map (
            O => \N__35501\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__7219\ : CascadeMux
    port map (
            O => \N__35498\,
            I => \N__35495\
        );

    \I__7218\ : InMux
    port map (
            O => \N__35495\,
            I => \N__35492\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__35492\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__7216\ : CascadeMux
    port map (
            O => \N__35489\,
            I => \N__35486\
        );

    \I__7215\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35483\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__35483\,
            I => \N__35480\
        );

    \I__7213\ : Odrv4
    port map (
            O => \N__35480\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__35477\,
            I => \N__35474\
        );

    \I__7211\ : InMux
    port map (
            O => \N__35474\,
            I => \N__35471\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__35471\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__7209\ : CascadeMux
    port map (
            O => \N__35468\,
            I => \N__35465\
        );

    \I__7208\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35462\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__35462\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__7206\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35456\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__35456\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__7204\ : InMux
    port map (
            O => \N__35453\,
            I => \N__35450\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__35450\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__7202\ : InMux
    port map (
            O => \N__35447\,
            I => \N__35443\
        );

    \I__7201\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35440\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__35443\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__35440\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__7198\ : CascadeMux
    port map (
            O => \N__35435\,
            I => \N__35432\
        );

    \I__7197\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__35429\,
            I => \N__35426\
        );

    \I__7195\ : Span4Mux_h
    port map (
            O => \N__35426\,
            I => \N__35422\
        );

    \I__7194\ : InMux
    port map (
            O => \N__35425\,
            I => \N__35419\
        );

    \I__7193\ : Odrv4
    port map (
            O => \N__35422\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__35419\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35414\,
            I => \N__35408\
        );

    \I__7190\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35408\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__35408\,
            I => \elapsed_time_ns_1_RNI2IIF91_0_28\
        );

    \I__7188\ : CascadeMux
    port map (
            O => \N__35405\,
            I => \N__35402\
        );

    \I__7187\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35399\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__35399\,
            I => \N__35395\
        );

    \I__7185\ : InMux
    port map (
            O => \N__35398\,
            I => \N__35392\
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__35395\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__35392\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35387\,
            I => \N__35383\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35386\,
            I => \N__35379\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__35383\,
            I => \N__35376\
        );

    \I__7179\ : InMux
    port map (
            O => \N__35382\,
            I => \N__35373\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__35379\,
            I => \N__35370\
        );

    \I__7177\ : Odrv4
    port map (
            O => \N__35376\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__35373\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__7175\ : Odrv4
    port map (
            O => \N__35370\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__7174\ : CascadeMux
    port map (
            O => \N__35363\,
            I => \N__35360\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35360\,
            I => \N__35357\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__35357\,
            I => \N__35353\
        );

    \I__7171\ : InMux
    port map (
            O => \N__35356\,
            I => \N__35350\
        );

    \I__7170\ : Span4Mux_v
    port map (
            O => \N__35353\,
            I => \N__35347\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__35350\,
            I => \N__35344\
        );

    \I__7168\ : Odrv4
    port map (
            O => \N__35347\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__7167\ : Odrv4
    port map (
            O => \N__35344\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35336\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35336\,
            I => \N__35332\
        );

    \I__7164\ : CascadeMux
    port map (
            O => \N__35335\,
            I => \N__35329\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__35332\,
            I => \N__35326\
        );

    \I__7162\ : InMux
    port map (
            O => \N__35329\,
            I => \N__35323\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__35326\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__35323\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__7159\ : CascadeMux
    port map (
            O => \N__35318\,
            I => \N__35315\
        );

    \I__7158\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35312\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35312\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__7156\ : CascadeMux
    port map (
            O => \N__35309\,
            I => \N__35306\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35303\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__35303\,
            I => \N__35300\
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__35300\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__7152\ : CascadeMux
    port map (
            O => \N__35297\,
            I => \N__35294\
        );

    \I__7151\ : InMux
    port map (
            O => \N__35294\,
            I => \N__35291\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35291\,
            I => \N__35288\
        );

    \I__7149\ : Odrv4
    port map (
            O => \N__35288\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35285\,
            I => \N__35282\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__35282\,
            I => \N__35279\
        );

    \I__7146\ : Span4Mux_v
    port map (
            O => \N__35279\,
            I => \N__35275\
        );

    \I__7145\ : InMux
    port map (
            O => \N__35278\,
            I => \N__35272\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__35275\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__35272\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__7142\ : CascadeMux
    port map (
            O => \N__35267\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35264\,
            I => \N__35261\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__35261\,
            I => \N__35258\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__35258\,
            I => \N__35254\
        );

    \I__7138\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35251\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__35254\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__35251\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__7135\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35243\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__35243\,
            I => \N__35240\
        );

    \I__7133\ : Span4Mux_h
    port map (
            O => \N__35240\,
            I => \N__35236\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35233\
        );

    \I__7131\ : Odrv4
    port map (
            O => \N__35236\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35233\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__7129\ : InMux
    port map (
            O => \N__35228\,
            I => \N__35225\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__35225\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35222\,
            I => \N__35218\
        );

    \I__7126\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35215\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__35218\,
            I => \elapsed_time_ns_1_RNI1HIF91_0_27\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__35215\,
            I => \elapsed_time_ns_1_RNI1HIF91_0_27\
        );

    \I__7123\ : CascadeMux
    port map (
            O => \N__35210\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\
        );

    \I__7122\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35204\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__35204\,
            I => \N__35201\
        );

    \I__7120\ : Span4Mux_h
    port map (
            O => \N__35201\,
            I => \N__35197\
        );

    \I__7119\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35194\
        );

    \I__7118\ : Span4Mux_v
    port map (
            O => \N__35197\,
            I => \N__35189\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35194\,
            I => \N__35186\
        );

    \I__7116\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35181\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35192\,
            I => \N__35181\
        );

    \I__7114\ : Odrv4
    port map (
            O => \N__35189\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__35186\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__35181\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__7111\ : InMux
    port map (
            O => \N__35174\,
            I => \N__35171\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35171\,
            I => \N__35168\
        );

    \I__7109\ : Span4Mux_h
    port map (
            O => \N__35168\,
            I => \N__35165\
        );

    \I__7108\ : Span4Mux_v
    port map (
            O => \N__35165\,
            I => \N__35161\
        );

    \I__7107\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35158\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__35161\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__35158\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__7104\ : CascadeMux
    port map (
            O => \N__35153\,
            I => \N__35150\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35147\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__35147\,
            I => \N__35143\
        );

    \I__7101\ : InMux
    port map (
            O => \N__35146\,
            I => \N__35140\
        );

    \I__7100\ : Odrv12
    port map (
            O => \N__35143\,
            I => \delay_measurement_inst.delay_tr_timer.N_381\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__35140\,
            I => \delay_measurement_inst.delay_tr_timer.N_381\
        );

    \I__7098\ : InMux
    port map (
            O => \N__35135\,
            I => \N__35132\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__35132\,
            I => \delay_measurement_inst.delay_tr_timer.N_358\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__35129\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\
        );

    \I__7095\ : InMux
    port map (
            O => \N__35126\,
            I => \N__35123\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__35123\,
            I => \N__35120\
        );

    \I__7093\ : Span4Mux_v
    port map (
            O => \N__35120\,
            I => \N__35116\
        );

    \I__7092\ : InMux
    port map (
            O => \N__35119\,
            I => \N__35113\
        );

    \I__7091\ : Odrv4
    port map (
            O => \N__35116\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__35113\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__7089\ : InMux
    port map (
            O => \N__35108\,
            I => \N__35104\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__35107\,
            I => \N__35100\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__35104\,
            I => \N__35097\
        );

    \I__7086\ : InMux
    port map (
            O => \N__35103\,
            I => \N__35094\
        );

    \I__7085\ : InMux
    port map (
            O => \N__35100\,
            I => \N__35091\
        );

    \I__7084\ : Span4Mux_h
    port map (
            O => \N__35097\,
            I => \N__35088\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__35094\,
            I => \N__35083\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__35091\,
            I => \N__35083\
        );

    \I__7081\ : Odrv4
    port map (
            O => \N__35088\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__7080\ : Odrv4
    port map (
            O => \N__35083\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__7079\ : CascadeMux
    port map (
            O => \N__35078\,
            I => \elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_\
        );

    \I__7078\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35072\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__35072\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35069\,
            I => \bfn_14_21_0_\
        );

    \I__7075\ : InMux
    port map (
            O => \N__35066\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__7074\ : CascadeMux
    port map (
            O => \N__35063\,
            I => \N__35060\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35060\,
            I => \N__35057\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__35057\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__7071\ : InMux
    port map (
            O => \N__35054\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__7070\ : InMux
    port map (
            O => \N__35051\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__7069\ : CascadeMux
    port map (
            O => \N__35048\,
            I => \N__35045\
        );

    \I__7068\ : InMux
    port map (
            O => \N__35045\,
            I => \N__35042\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__35042\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__7066\ : InMux
    port map (
            O => \N__35039\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__7065\ : InMux
    port map (
            O => \N__35036\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__7064\ : InMux
    port map (
            O => \N__35033\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__7063\ : InMux
    port map (
            O => \N__35030\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35027\,
            I => \N__35024\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__35024\,
            I => \N__35021\
        );

    \I__7060\ : Odrv12
    port map (
            O => \N__35021\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__35018\,
            I => \N__35015\
        );

    \I__7058\ : InMux
    port map (
            O => \N__35015\,
            I => \N__35012\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__35012\,
            I => \N__35009\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__35009\,
            I => \N__35006\
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__35006\,
            I => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\
        );

    \I__7054\ : InMux
    port map (
            O => \N__35003\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__7053\ : CascadeMux
    port map (
            O => \N__35000\,
            I => \N__34997\
        );

    \I__7052\ : InMux
    port map (
            O => \N__34997\,
            I => \N__34994\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__34994\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__7050\ : InMux
    port map (
            O => \N__34991\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__7049\ : InMux
    port map (
            O => \N__34988\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__7048\ : InMux
    port map (
            O => \N__34985\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__7047\ : InMux
    port map (
            O => \N__34982\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__7046\ : InMux
    port map (
            O => \N__34979\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__7045\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34973\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__34973\,
            I => \N__34970\
        );

    \I__7043\ : Odrv4
    port map (
            O => \N__34970\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__7042\ : InMux
    port map (
            O => \N__34967\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__7041\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34960\
        );

    \I__7040\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34957\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__34960\,
            I => \N__34954\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__34957\,
            I => \N__34951\
        );

    \I__7037\ : Odrv4
    port map (
            O => \N__34954\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__7036\ : Odrv4
    port map (
            O => \N__34951\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__7035\ : InMux
    port map (
            O => \N__34946\,
            I => \N__34943\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__34943\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__7033\ : InMux
    port map (
            O => \N__34940\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__7032\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34934\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__34934\,
            I => \N__34931\
        );

    \I__7030\ : Odrv4
    port map (
            O => \N__34931\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__7029\ : InMux
    port map (
            O => \N__34928\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__7028\ : InMux
    port map (
            O => \N__34925\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__7027\ : InMux
    port map (
            O => \N__34922\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__7026\ : InMux
    port map (
            O => \N__34919\,
            I => \bfn_14_17_0_\
        );

    \I__7025\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34913\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__34913\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__7023\ : InMux
    port map (
            O => \N__34910\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__7022\ : InMux
    port map (
            O => \N__34907\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__7021\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34901\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__34901\,
            I => \N__34898\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__34898\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__7018\ : InMux
    port map (
            O => \N__34895\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__34892\,
            I => \N__34889\
        );

    \I__7016\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34886\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__34886\,
            I => \N__34883\
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__34883\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__7013\ : InMux
    port map (
            O => \N__34880\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__7012\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34874\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__34874\,
            I => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\
        );

    \I__7010\ : InMux
    port map (
            O => \N__34871\,
            I => \N__34868\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__34868\,
            I => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\
        );

    \I__7008\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34862\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__34862\,
            I => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\
        );

    \I__7006\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34856\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__34856\,
            I => \N__34853\
        );

    \I__7004\ : Odrv4
    port map (
            O => \N__34853\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__34850\,
            I => \N__34847\
        );

    \I__7002\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34844\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__34844\,
            I => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\
        );

    \I__7000\ : CascadeMux
    port map (
            O => \N__34841\,
            I => \N__34838\
        );

    \I__6999\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34835\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__34835\,
            I => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\
        );

    \I__6997\ : CascadeMux
    port map (
            O => \N__34832\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_\
        );

    \I__6996\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34822\
        );

    \I__6995\ : InMux
    port map (
            O => \N__34828\,
            I => \N__34822\
        );

    \I__6994\ : InMux
    port map (
            O => \N__34827\,
            I => \N__34819\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__34822\,
            I => \N__34816\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__34819\,
            I => \N__34813\
        );

    \I__6991\ : Span4Mux_h
    port map (
            O => \N__34816\,
            I => \N__34809\
        );

    \I__6990\ : Span4Mux_v
    port map (
            O => \N__34813\,
            I => \N__34806\
        );

    \I__6989\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34803\
        );

    \I__6988\ : Span4Mux_v
    port map (
            O => \N__34809\,
            I => \N__34798\
        );

    \I__6987\ : Span4Mux_h
    port map (
            O => \N__34806\,
            I => \N__34793\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__34803\,
            I => \N__34793\
        );

    \I__6985\ : InMux
    port map (
            O => \N__34802\,
            I => \N__34790\
        );

    \I__6984\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34787\
        );

    \I__6983\ : Odrv4
    port map (
            O => \N__34798\,
            I => phase_controller_inst1_state_4
        );

    \I__6982\ : Odrv4
    port map (
            O => \N__34793\,
            I => phase_controller_inst1_state_4
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__34790\,
            I => phase_controller_inst1_state_4
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__34787\,
            I => phase_controller_inst1_state_4
        );

    \I__6979\ : CascadeMux
    port map (
            O => \N__34778\,
            I => \N__34775\
        );

    \I__6978\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34772\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__34772\,
            I => \phase_controller_inst2.stoper_tr.un1_start_latched2_0\
        );

    \I__6976\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34765\
        );

    \I__6975\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34762\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34756\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__34762\,
            I => \N__34756\
        );

    \I__6972\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34753\
        );

    \I__6971\ : Span4Mux_v
    port map (
            O => \N__34756\,
            I => \N__34750\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__34753\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6969\ : Odrv4
    port map (
            O => \N__34750\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6968\ : CascadeMux
    port map (
            O => \N__34745\,
            I => \N__34742\
        );

    \I__6967\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34739\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__34739\,
            I => \phase_controller_inst2.stoper_tr.running_1_sqmuxa\
        );

    \I__6965\ : InMux
    port map (
            O => \N__34736\,
            I => \N__34731\
        );

    \I__6964\ : InMux
    port map (
            O => \N__34735\,
            I => \N__34726\
        );

    \I__6963\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34726\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__34731\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__34726\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__6960\ : InMux
    port map (
            O => \N__34721\,
            I => \N__34709\
        );

    \I__6959\ : InMux
    port map (
            O => \N__34720\,
            I => \N__34709\
        );

    \I__6958\ : InMux
    port map (
            O => \N__34719\,
            I => \N__34709\
        );

    \I__6957\ : InMux
    port map (
            O => \N__34718\,
            I => \N__34702\
        );

    \I__6956\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34702\
        );

    \I__6955\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34702\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__34709\,
            I => \N__34697\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__34702\,
            I => \N__34697\
        );

    \I__6952\ : Span4Mux_h
    port map (
            O => \N__34697\,
            I => \N__34693\
        );

    \I__6951\ : InMux
    port map (
            O => \N__34696\,
            I => \N__34690\
        );

    \I__6950\ : Span4Mux_v
    port map (
            O => \N__34693\,
            I => \N__34687\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__34690\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__34687\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__6947\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34672\
        );

    \I__6946\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34672\
        );

    \I__6945\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34669\
        );

    \I__6944\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34664\
        );

    \I__6943\ : InMux
    port map (
            O => \N__34678\,
            I => \N__34664\
        );

    \I__6942\ : CascadeMux
    port map (
            O => \N__34677\,
            I => \N__34661\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__34672\,
            I => \N__34657\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__34669\,
            I => \N__34651\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__34664\,
            I => \N__34651\
        );

    \I__6938\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34646\
        );

    \I__6937\ : InMux
    port map (
            O => \N__34660\,
            I => \N__34646\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__34657\,
            I => \N__34643\
        );

    \I__6935\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34640\
        );

    \I__6934\ : Span4Mux_v
    port map (
            O => \N__34651\,
            I => \N__34637\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__34646\,
            I => \N__34632\
        );

    \I__6932\ : Span4Mux_v
    port map (
            O => \N__34643\,
            I => \N__34632\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__34640\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__34637\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__34632\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__6928\ : InMux
    port map (
            O => \N__34625\,
            I => \N__34622\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__34622\,
            I => \N__34619\
        );

    \I__6926\ : Span4Mux_v
    port map (
            O => \N__34619\,
            I => \N__34616\
        );

    \I__6925\ : Span4Mux_h
    port map (
            O => \N__34616\,
            I => \N__34613\
        );

    \I__6924\ : Span4Mux_h
    port map (
            O => \N__34613\,
            I => \N__34609\
        );

    \I__6923\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34606\
        );

    \I__6922\ : Odrv4
    port map (
            O => \N__34609\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__34606\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__34601\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__6919\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34595\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__34595\,
            I => \N__34592\
        );

    \I__6917\ : Span4Mux_v
    port map (
            O => \N__34592\,
            I => \N__34589\
        );

    \I__6916\ : Span4Mux_h
    port map (
            O => \N__34589\,
            I => \N__34586\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__34586\,
            I => \N__34581\
        );

    \I__6914\ : InMux
    port map (
            O => \N__34585\,
            I => \N__34576\
        );

    \I__6913\ : InMux
    port map (
            O => \N__34584\,
            I => \N__34576\
        );

    \I__6912\ : Odrv4
    port map (
            O => \N__34581\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__34576\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__6910\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34568\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__34568\,
            I => \N__34565\
        );

    \I__6908\ : Odrv12
    port map (
            O => \N__34565\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__34562\,
            I => \N__34558\
        );

    \I__6906\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34555\
        );

    \I__6905\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34552\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__34555\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__34552\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__34547\,
            I => \N__34544\
        );

    \I__6901\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34541\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__34541\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23\
        );

    \I__6899\ : CascadeMux
    port map (
            O => \N__34538\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34535\,
            I => \N__34531\
        );

    \I__6897\ : InMux
    port map (
            O => \N__34534\,
            I => \N__34528\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__34531\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34528\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__6894\ : InMux
    port map (
            O => \N__34523\,
            I => \N__34520\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__34520\,
            I => \N__34517\
        );

    \I__6892\ : Odrv4
    port map (
            O => \N__34517\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__6891\ : CascadeMux
    port map (
            O => \N__34514\,
            I => \phase_controller_inst1.N_55_cascade_\
        );

    \I__6890\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34502\
        );

    \I__6889\ : InMux
    port map (
            O => \N__34510\,
            I => \N__34502\
        );

    \I__6888\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34502\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__34502\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6886\ : CascadeMux
    port map (
            O => \N__34499\,
            I => \N__34495\
        );

    \I__6885\ : InMux
    port map (
            O => \N__34498\,
            I => \N__34490\
        );

    \I__6884\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34490\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__34490\,
            I => \N__34487\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__34487\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__6881\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34478\
        );

    \I__6880\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34478\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34478\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__6878\ : InMux
    port map (
            O => \N__34475\,
            I => \N__34468\
        );

    \I__6877\ : InMux
    port map (
            O => \N__34474\,
            I => \N__34468\
        );

    \I__6876\ : InMux
    port map (
            O => \N__34473\,
            I => \N__34465\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__34468\,
            I => \N__34462\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__34465\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\
        );

    \I__6873\ : Odrv4
    port map (
            O => \N__34462\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\
        );

    \I__6872\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34454\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__34454\,
            I => \delay_measurement_inst.delay_tr_timer.N_347\
        );

    \I__6870\ : CascadeMux
    port map (
            O => \N__34451\,
            I => \delay_measurement_inst.delay_tr_timer.N_347_cascade_\
        );

    \I__6869\ : CascadeMux
    port map (
            O => \N__34448\,
            I => \N__34443\
        );

    \I__6868\ : InMux
    port map (
            O => \N__34447\,
            I => \N__34440\
        );

    \I__6867\ : InMux
    port map (
            O => \N__34446\,
            I => \N__34435\
        );

    \I__6866\ : InMux
    port map (
            O => \N__34443\,
            I => \N__34435\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__34440\,
            I => \N__34432\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__34435\,
            I => \N__34429\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__34432\,
            I => \delay_measurement_inst.delay_tr_timer.N_365\
        );

    \I__6862\ : Odrv12
    port map (
            O => \N__34429\,
            I => \delay_measurement_inst.delay_tr_timer.N_365\
        );

    \I__6861\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34420\
        );

    \I__6860\ : CascadeMux
    port map (
            O => \N__34423\,
            I => \N__34417\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__34420\,
            I => \N__34414\
        );

    \I__6858\ : InMux
    port map (
            O => \N__34417\,
            I => \N__34411\
        );

    \I__6857\ : Odrv4
    port map (
            O => \N__34414\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__34411\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__6855\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34401\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34405\,
            I => \N__34396\
        );

    \I__6853\ : InMux
    port map (
            O => \N__34404\,
            I => \N__34396\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__34401\,
            I => \N__34393\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__34396\,
            I => \N__34390\
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__34393\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\
        );

    \I__6849\ : Odrv12
    port map (
            O => \N__34390\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\
        );

    \I__6848\ : InMux
    port map (
            O => \N__34385\,
            I => \N__34381\
        );

    \I__6847\ : InMux
    port map (
            O => \N__34384\,
            I => \N__34378\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__34381\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__34378\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34373\,
            I => \N__34370\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34370\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6\
        );

    \I__6842\ : CascadeMux
    port map (
            O => \N__34367\,
            I => \N__34363\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34360\
        );

    \I__6840\ : InMux
    port map (
            O => \N__34363\,
            I => \N__34357\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__34360\,
            I => \delay_measurement_inst.delay_tr_timer.N_341\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__34357\,
            I => \delay_measurement_inst.delay_tr_timer.N_341\
        );

    \I__6837\ : CascadeMux
    port map (
            O => \N__34352\,
            I => \N__34348\
        );

    \I__6836\ : InMux
    port map (
            O => \N__34351\,
            I => \N__34345\
        );

    \I__6835\ : InMux
    port map (
            O => \N__34348\,
            I => \N__34342\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34345\,
            I => \N__34339\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__34342\,
            I => \N__34335\
        );

    \I__6832\ : Span4Mux_v
    port map (
            O => \N__34339\,
            I => \N__34332\
        );

    \I__6831\ : InMux
    port map (
            O => \N__34338\,
            I => \N__34329\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__34335\,
            I => \N__34326\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__34332\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__34329\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__34326\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__6826\ : InMux
    port map (
            O => \N__34319\,
            I => \N__34312\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34312\
        );

    \I__6824\ : InMux
    port map (
            O => \N__34317\,
            I => \N__34309\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__34312\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__34309\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__6821\ : CEMux
    port map (
            O => \N__34304\,
            I => \N__34286\
        );

    \I__6820\ : CEMux
    port map (
            O => \N__34303\,
            I => \N__34286\
        );

    \I__6819\ : CEMux
    port map (
            O => \N__34302\,
            I => \N__34286\
        );

    \I__6818\ : CEMux
    port map (
            O => \N__34301\,
            I => \N__34286\
        );

    \I__6817\ : CEMux
    port map (
            O => \N__34300\,
            I => \N__34286\
        );

    \I__6816\ : CEMux
    port map (
            O => \N__34299\,
            I => \N__34286\
        );

    \I__6815\ : GlobalMux
    port map (
            O => \N__34286\,
            I => \N__34283\
        );

    \I__6814\ : gio2CtrlBuf
    port map (
            O => \N__34283\,
            I => \delay_measurement_inst.delay_tr_timer.N_434_i_g\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34277\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34274\
        );

    \I__6811\ : Odrv4
    port map (
            O => \N__34274\,
            I => \delay_measurement_inst.delay_tr_timer.N_348\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34271\,
            I => \N__34267\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34264\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__34267\,
            I => \delay_measurement_inst.delay_tr_timer.N_367\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__34264\,
            I => \delay_measurement_inst.delay_tr_timer.N_367\
        );

    \I__6806\ : CascadeMux
    port map (
            O => \N__34259\,
            I => \delay_measurement_inst.delay_tr_timer.N_349_cascade_\
        );

    \I__6805\ : CascadeMux
    port map (
            O => \N__34256\,
            I => \delay_measurement_inst.delay_tr_timer.N_363_cascade_\
        );

    \I__6804\ : CascadeMux
    port map (
            O => \N__34253\,
            I => \N__34249\
        );

    \I__6803\ : InMux
    port map (
            O => \N__34252\,
            I => \N__34246\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34243\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__34246\,
            I => \delay_measurement_inst.delay_tr_timer.N_380\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__34243\,
            I => \delay_measurement_inst.delay_tr_timer.N_380\
        );

    \I__6799\ : CascadeMux
    port map (
            O => \N__34238\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_\
        );

    \I__6798\ : CascadeMux
    port map (
            O => \N__34235\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_\
        );

    \I__6797\ : InMux
    port map (
            O => \N__34232\,
            I => \N__34225\
        );

    \I__6796\ : InMux
    port map (
            O => \N__34231\,
            I => \N__34225\
        );

    \I__6795\ : InMux
    port map (
            O => \N__34230\,
            I => \N__34222\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34225\,
            I => \delay_measurement_inst.delay_tr_timer.N_378\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__34222\,
            I => \delay_measurement_inst.delay_tr_timer.N_378\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34217\,
            I => \N__34214\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34214\,
            I => \N__34211\
        );

    \I__6790\ : Odrv4
    port map (
            O => \N__34211\,
            I => \delay_measurement_inst.delay_tr_timer.N_359_1\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34202\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34202\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34202\,
            I => \N__34198\
        );

    \I__6786\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34195\
        );

    \I__6785\ : Span4Mux_v
    port map (
            O => \N__34198\,
            I => \N__34192\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__34195\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__6783\ : Odrv4
    port map (
            O => \N__34192\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__34187\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\
        );

    \I__6781\ : CascadeMux
    port map (
            O => \N__34184\,
            I => \delay_measurement_inst.delay_tr_timer.N_359_1_cascade_\
        );

    \I__6780\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34178\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__34178\,
            I => \delay_measurement_inst.delay_tr_timer.N_345\
        );

    \I__6778\ : CascadeMux
    port map (
            O => \N__34175\,
            I => \delay_measurement_inst.delay_tr_timer.N_345_cascade_\
        );

    \I__6777\ : CascadeMux
    port map (
            O => \N__34172\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\
        );

    \I__6776\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34166\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__34166\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\
        );

    \I__6774\ : InMux
    port map (
            O => \N__34163\,
            I => \N__34160\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__34160\,
            I => \N__34156\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34153\
        );

    \I__6771\ : Span4Mux_s1_v
    port map (
            O => \N__34156\,
            I => \N__34148\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__34153\,
            I => \N__34148\
        );

    \I__6769\ : Span4Mux_v
    port map (
            O => \N__34148\,
            I => \N__34143\
        );

    \I__6768\ : InMux
    port map (
            O => \N__34147\,
            I => \N__34140\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34146\,
            I => \N__34137\
        );

    \I__6766\ : Span4Mux_h
    port map (
            O => \N__34143\,
            I => \N__34134\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__34140\,
            I => \N__34131\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__34137\,
            I => \N__34128\
        );

    \I__6763\ : Sp12to4
    port map (
            O => \N__34134\,
            I => \N__34125\
        );

    \I__6762\ : Span4Mux_v
    port map (
            O => \N__34131\,
            I => \N__34122\
        );

    \I__6761\ : Span4Mux_v
    port map (
            O => \N__34128\,
            I => \N__34119\
        );

    \I__6760\ : Span12Mux_v
    port map (
            O => \N__34125\,
            I => \N__34116\
        );

    \I__6759\ : Sp12to4
    port map (
            O => \N__34122\,
            I => \N__34113\
        );

    \I__6758\ : Span4Mux_h
    port map (
            O => \N__34119\,
            I => \N__34110\
        );

    \I__6757\ : Span12Mux_v
    port map (
            O => \N__34116\,
            I => \N__34107\
        );

    \I__6756\ : Span12Mux_h
    port map (
            O => \N__34113\,
            I => \N__34102\
        );

    \I__6755\ : Sp12to4
    port map (
            O => \N__34110\,
            I => \N__34102\
        );

    \I__6754\ : Span12Mux_h
    port map (
            O => \N__34107\,
            I => \N__34099\
        );

    \I__6753\ : Span12Mux_v
    port map (
            O => \N__34102\,
            I => \N__34096\
        );

    \I__6752\ : Odrv12
    port map (
            O => \N__34099\,
            I => start_stop_c
        );

    \I__6751\ : Odrv12
    port map (
            O => \N__34096\,
            I => start_stop_c
        );

    \I__6750\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34088\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__34088\,
            I => \N__34085\
        );

    \I__6748\ : Span4Mux_v
    port map (
            O => \N__34085\,
            I => \N__34082\
        );

    \I__6747\ : Span4Mux_v
    port map (
            O => \N__34082\,
            I => \N__34079\
        );

    \I__6746\ : Odrv4
    port map (
            O => \N__34079\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__6745\ : IoInMux
    port map (
            O => \N__34076\,
            I => \N__34073\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__34073\,
            I => \N__34070\
        );

    \I__6743\ : Span4Mux_s2_v
    port map (
            O => \N__34070\,
            I => \N__34067\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__34067\,
            I => s2_phy_c
        );

    \I__6741\ : InMux
    port map (
            O => \N__34064\,
            I => \N__34060\
        );

    \I__6740\ : InMux
    port map (
            O => \N__34063\,
            I => \N__34056\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__34060\,
            I => \N__34053\
        );

    \I__6738\ : InMux
    port map (
            O => \N__34059\,
            I => \N__34050\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__34056\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__6736\ : Odrv12
    port map (
            O => \N__34053\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__34050\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__6734\ : InMux
    port map (
            O => \N__34043\,
            I => \N__34040\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__34040\,
            I => \N__34037\
        );

    \I__6732\ : Span4Mux_h
    port map (
            O => \N__34037\,
            I => \N__34033\
        );

    \I__6731\ : InMux
    port map (
            O => \N__34036\,
            I => \N__34030\
        );

    \I__6730\ : Span4Mux_v
    port map (
            O => \N__34033\,
            I => \N__34021\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__34030\,
            I => \N__34021\
        );

    \I__6728\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34018\
        );

    \I__6727\ : InMux
    port map (
            O => \N__34028\,
            I => \N__34013\
        );

    \I__6726\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34013\
        );

    \I__6725\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34010\
        );

    \I__6724\ : Odrv4
    port map (
            O => \N__34021\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__34018\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__34013\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__34010\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6720\ : CascadeMux
    port map (
            O => \N__34001\,
            I => \N__33997\
        );

    \I__6719\ : InMux
    port map (
            O => \N__34000\,
            I => \N__33993\
        );

    \I__6718\ : InMux
    port map (
            O => \N__33997\,
            I => \N__33988\
        );

    \I__6717\ : InMux
    port map (
            O => \N__33996\,
            I => \N__33988\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__33993\,
            I => \N__33985\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__33988\,
            I => \N__33982\
        );

    \I__6714\ : Sp12to4
    port map (
            O => \N__33985\,
            I => \N__33979\
        );

    \I__6713\ : Span4Mux_v
    port map (
            O => \N__33982\,
            I => \N__33976\
        );

    \I__6712\ : Span12Mux_h
    port map (
            O => \N__33979\,
            I => \N__33973\
        );

    \I__6711\ : Span4Mux_v
    port map (
            O => \N__33976\,
            I => \N__33970\
        );

    \I__6710\ : Span12Mux_v
    port map (
            O => \N__33973\,
            I => \N__33967\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__33970\,
            I => \il_min_comp2_D2\
        );

    \I__6708\ : Odrv12
    port map (
            O => \N__33967\,
            I => \il_min_comp2_D2\
        );

    \I__6707\ : InMux
    port map (
            O => \N__33962\,
            I => \N__33959\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__33959\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa\
        );

    \I__6705\ : CascadeMux
    port map (
            O => \N__33956\,
            I => \N__33953\
        );

    \I__6704\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33950\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__33950\,
            I => \N__33947\
        );

    \I__6702\ : Sp12to4
    port map (
            O => \N__33947\,
            I => \N__33944\
        );

    \I__6701\ : Odrv12
    port map (
            O => \N__33944\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__6700\ : CascadeMux
    port map (
            O => \N__33941\,
            I => \N__33936\
        );

    \I__6699\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33933\
        );

    \I__6698\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33930\
        );

    \I__6697\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33926\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__33933\,
            I => \N__33923\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__33930\,
            I => \N__33920\
        );

    \I__6694\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33917\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__33926\,
            I => \N__33914\
        );

    \I__6692\ : Span4Mux_v
    port map (
            O => \N__33923\,
            I => \N__33905\
        );

    \I__6691\ : Span4Mux_v
    port map (
            O => \N__33920\,
            I => \N__33905\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__33917\,
            I => \N__33905\
        );

    \I__6689\ : Span4Mux_v
    port map (
            O => \N__33914\,
            I => \N__33905\
        );

    \I__6688\ : Odrv4
    port map (
            O => \N__33905\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16\
        );

    \I__6687\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33899\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33895\
        );

    \I__6685\ : CascadeMux
    port map (
            O => \N__33898\,
            I => \N__33892\
        );

    \I__6684\ : Span4Mux_h
    port map (
            O => \N__33895\,
            I => \N__33888\
        );

    \I__6683\ : InMux
    port map (
            O => \N__33892\,
            I => \N__33883\
        );

    \I__6682\ : InMux
    port map (
            O => \N__33891\,
            I => \N__33883\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__33888\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__33883\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__6679\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33875\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__33875\,
            I => \N__33872\
        );

    \I__6677\ : Span4Mux_h
    port map (
            O => \N__33872\,
            I => \N__33869\
        );

    \I__6676\ : Odrv4
    port map (
            O => \N__33869\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16\
        );

    \I__6675\ : CascadeMux
    port map (
            O => \N__33866\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__6674\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33860\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__33860\,
            I => \N__33857\
        );

    \I__6672\ : Span4Mux_v
    port map (
            O => \N__33857\,
            I => \N__33854\
        );

    \I__6671\ : Odrv4
    port map (
            O => \N__33854\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__6670\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33848\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__33848\,
            I => \N__33844\
        );

    \I__6668\ : InMux
    port map (
            O => \N__33847\,
            I => \N__33841\
        );

    \I__6667\ : Span4Mux_h
    port map (
            O => \N__33844\,
            I => \N__33837\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__33841\,
            I => \N__33834\
        );

    \I__6665\ : InMux
    port map (
            O => \N__33840\,
            I => \N__33831\
        );

    \I__6664\ : Span4Mux_v
    port map (
            O => \N__33837\,
            I => \N__33828\
        );

    \I__6663\ : Odrv4
    port map (
            O => \N__33834\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__33831\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__6661\ : Odrv4
    port map (
            O => \N__33828\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__6660\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33816\
        );

    \I__6659\ : InMux
    port map (
            O => \N__33820\,
            I => \N__33810\
        );

    \I__6658\ : InMux
    port map (
            O => \N__33819\,
            I => \N__33810\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__33816\,
            I => \N__33807\
        );

    \I__6656\ : InMux
    port map (
            O => \N__33815\,
            I => \N__33804\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__33810\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__6654\ : Odrv4
    port map (
            O => \N__33807\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__33804\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__6652\ : ClkMux
    port map (
            O => \N__33797\,
            I => \N__33794\
        );

    \I__6651\ : GlobalMux
    port map (
            O => \N__33794\,
            I => \N__33791\
        );

    \I__6650\ : gio2CtrlBuf
    port map (
            O => \N__33791\,
            I => delay_tr_input_c_g
        );

    \I__6649\ : InMux
    port map (
            O => \N__33788\,
            I => \N__33785\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__33785\,
            I => \N__33782\
        );

    \I__6647\ : Span4Mux_v
    port map (
            O => \N__33782\,
            I => \N__33779\
        );

    \I__6646\ : Odrv4
    port map (
            O => \N__33779\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__6645\ : CascadeMux
    port map (
            O => \N__33776\,
            I => \N__33770\
        );

    \I__6644\ : CascadeMux
    port map (
            O => \N__33775\,
            I => \N__33767\
        );

    \I__6643\ : InMux
    port map (
            O => \N__33774\,
            I => \N__33752\
        );

    \I__6642\ : InMux
    port map (
            O => \N__33773\,
            I => \N__33749\
        );

    \I__6641\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33746\
        );

    \I__6640\ : InMux
    port map (
            O => \N__33767\,
            I => \N__33738\
        );

    \I__6639\ : InMux
    port map (
            O => \N__33766\,
            I => \N__33735\
        );

    \I__6638\ : InMux
    port map (
            O => \N__33765\,
            I => \N__33728\
        );

    \I__6637\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33728\
        );

    \I__6636\ : InMux
    port map (
            O => \N__33763\,
            I => \N__33728\
        );

    \I__6635\ : CascadeMux
    port map (
            O => \N__33762\,
            I => \N__33722\
        );

    \I__6634\ : CascadeMux
    port map (
            O => \N__33761\,
            I => \N__33719\
        );

    \I__6633\ : CascadeMux
    port map (
            O => \N__33760\,
            I => \N__33713\
        );

    \I__6632\ : CascadeMux
    port map (
            O => \N__33759\,
            I => \N__33709\
        );

    \I__6631\ : CascadeMux
    port map (
            O => \N__33758\,
            I => \N__33704\
        );

    \I__6630\ : CascadeMux
    port map (
            O => \N__33757\,
            I => \N__33699\
        );

    \I__6629\ : CascadeMux
    port map (
            O => \N__33756\,
            I => \N__33696\
        );

    \I__6628\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33688\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__33752\,
            I => \N__33685\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__33749\,
            I => \N__33680\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__33746\,
            I => \N__33680\
        );

    \I__6624\ : CascadeMux
    port map (
            O => \N__33745\,
            I => \N__33673\
        );

    \I__6623\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33666\
        );

    \I__6622\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33661\
        );

    \I__6621\ : InMux
    port map (
            O => \N__33742\,
            I => \N__33661\
        );

    \I__6620\ : InMux
    port map (
            O => \N__33741\,
            I => \N__33658\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__33738\,
            I => \N__33651\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__33735\,
            I => \N__33651\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__33728\,
            I => \N__33651\
        );

    \I__6616\ : InMux
    port map (
            O => \N__33727\,
            I => \N__33644\
        );

    \I__6615\ : InMux
    port map (
            O => \N__33726\,
            I => \N__33644\
        );

    \I__6614\ : InMux
    port map (
            O => \N__33725\,
            I => \N__33644\
        );

    \I__6613\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33631\
        );

    \I__6612\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33631\
        );

    \I__6611\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33631\
        );

    \I__6610\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33631\
        );

    \I__6609\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33631\
        );

    \I__6608\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33631\
        );

    \I__6607\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33616\
        );

    \I__6606\ : InMux
    port map (
            O => \N__33709\,
            I => \N__33616\
        );

    \I__6605\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33616\
        );

    \I__6604\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33616\
        );

    \I__6603\ : InMux
    port map (
            O => \N__33704\,
            I => \N__33616\
        );

    \I__6602\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33616\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33702\,
            I => \N__33616\
        );

    \I__6600\ : InMux
    port map (
            O => \N__33699\,
            I => \N__33603\
        );

    \I__6599\ : InMux
    port map (
            O => \N__33696\,
            I => \N__33603\
        );

    \I__6598\ : InMux
    port map (
            O => \N__33695\,
            I => \N__33603\
        );

    \I__6597\ : InMux
    port map (
            O => \N__33694\,
            I => \N__33603\
        );

    \I__6596\ : InMux
    port map (
            O => \N__33693\,
            I => \N__33603\
        );

    \I__6595\ : InMux
    port map (
            O => \N__33692\,
            I => \N__33603\
        );

    \I__6594\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33594\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__33688\,
            I => \N__33587\
        );

    \I__6592\ : Span4Mux_v
    port map (
            O => \N__33685\,
            I => \N__33587\
        );

    \I__6591\ : Span4Mux_v
    port map (
            O => \N__33680\,
            I => \N__33587\
        );

    \I__6590\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33584\
        );

    \I__6589\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33579\
        );

    \I__6588\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33579\
        );

    \I__6587\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33566\
        );

    \I__6586\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33566\
        );

    \I__6585\ : InMux
    port map (
            O => \N__33672\,
            I => \N__33566\
        );

    \I__6584\ : InMux
    port map (
            O => \N__33671\,
            I => \N__33566\
        );

    \I__6583\ : InMux
    port map (
            O => \N__33670\,
            I => \N__33566\
        );

    \I__6582\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33566\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__33666\,
            I => \N__33561\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__33661\,
            I => \N__33561\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__33658\,
            I => \N__33548\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__33651\,
            I => \N__33548\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__33644\,
            I => \N__33548\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__33631\,
            I => \N__33548\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__33616\,
            I => \N__33548\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__33603\,
            I => \N__33548\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33545\
        );

    \I__6572\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33534\
        );

    \I__6571\ : InMux
    port map (
            O => \N__33600\,
            I => \N__33534\
        );

    \I__6570\ : InMux
    port map (
            O => \N__33599\,
            I => \N__33534\
        );

    \I__6569\ : InMux
    port map (
            O => \N__33598\,
            I => \N__33534\
        );

    \I__6568\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33534\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__33594\,
            I => \N__33529\
        );

    \I__6566\ : Span4Mux_h
    port map (
            O => \N__33587\,
            I => \N__33529\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__33584\,
            I => \N__33526\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__33579\,
            I => \N__33523\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__33566\,
            I => \N__33516\
        );

    \I__6562\ : Span4Mux_v
    port map (
            O => \N__33561\,
            I => \N__33516\
        );

    \I__6561\ : Span4Mux_v
    port map (
            O => \N__33548\,
            I => \N__33516\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__33545\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__33534\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6558\ : Odrv4
    port map (
            O => \N__33529\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6557\ : Odrv4
    port map (
            O => \N__33526\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6556\ : Odrv12
    port map (
            O => \N__33523\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6555\ : Odrv4
    port map (
            O => \N__33516\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__33503\,
            I => \N__33498\
        );

    \I__6553\ : InMux
    port map (
            O => \N__33502\,
            I => \N__33495\
        );

    \I__6552\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33490\
        );

    \I__6551\ : InMux
    port map (
            O => \N__33498\,
            I => \N__33490\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__33495\,
            I => \N__33485\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__33490\,
            I => \N__33485\
        );

    \I__6548\ : Span4Mux_h
    port map (
            O => \N__33485\,
            I => \N__33482\
        );

    \I__6547\ : Span4Mux_h
    port map (
            O => \N__33482\,
            I => \N__33479\
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__33479\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_0_12\
        );

    \I__6545\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33473\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__33473\,
            I => \N__33470\
        );

    \I__6543\ : Span4Mux_h
    port map (
            O => \N__33470\,
            I => \N__33467\
        );

    \I__6542\ : Odrv4
    port map (
            O => \N__33467\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__6541\ : InMux
    port map (
            O => \N__33464\,
            I => \N__33457\
        );

    \I__6540\ : InMux
    port map (
            O => \N__33463\,
            I => \N__33457\
        );

    \I__6539\ : InMux
    port map (
            O => \N__33462\,
            I => \N__33454\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__33457\,
            I => \N__33451\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__33454\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__6536\ : Odrv12
    port map (
            O => \N__33451\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__33446\,
            I => \N__33443\
        );

    \I__6534\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33439\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33442\,
            I => \N__33436\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__33439\,
            I => \N__33433\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__33436\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__6530\ : Odrv12
    port map (
            O => \N__33433\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__6529\ : InMux
    port map (
            O => \N__33428\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__6528\ : InMux
    port map (
            O => \N__33425\,
            I => \N__33421\
        );

    \I__6527\ : InMux
    port map (
            O => \N__33424\,
            I => \N__33418\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__33421\,
            I => \N__33415\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__33418\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__6524\ : Odrv12
    port map (
            O => \N__33415\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__6523\ : CascadeMux
    port map (
            O => \N__33410\,
            I => \N__33407\
        );

    \I__6522\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33403\
        );

    \I__6521\ : InMux
    port map (
            O => \N__33406\,
            I => \N__33400\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__33403\,
            I => \N__33394\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__33400\,
            I => \N__33394\
        );

    \I__6518\ : InMux
    port map (
            O => \N__33399\,
            I => \N__33391\
        );

    \I__6517\ : Span4Mux_v
    port map (
            O => \N__33394\,
            I => \N__33388\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__33391\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__6515\ : Odrv4
    port map (
            O => \N__33388\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__6514\ : InMux
    port map (
            O => \N__33383\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__6513\ : InMux
    port map (
            O => \N__33380\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__6512\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33373\
        );

    \I__6511\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33370\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__33373\,
            I => \N__33367\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__33370\,
            I => \N__33361\
        );

    \I__6508\ : Span4Mux_h
    port map (
            O => \N__33367\,
            I => \N__33361\
        );

    \I__6507\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33357\
        );

    \I__6506\ : Span4Mux_v
    port map (
            O => \N__33361\,
            I => \N__33354\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33360\,
            I => \N__33351\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__33357\,
            I => \N__33348\
        );

    \I__6503\ : Span4Mux_v
    port map (
            O => \N__33354\,
            I => \N__33345\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__33351\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6501\ : Odrv4
    port map (
            O => \N__33348\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6500\ : Odrv4
    port map (
            O => \N__33345\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6499\ : CEMux
    port map (
            O => \N__33338\,
            I => \N__33332\
        );

    \I__6498\ : CEMux
    port map (
            O => \N__33337\,
            I => \N__33329\
        );

    \I__6497\ : CEMux
    port map (
            O => \N__33336\,
            I => \N__33326\
        );

    \I__6496\ : CEMux
    port map (
            O => \N__33335\,
            I => \N__33323\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__33332\,
            I => \N__33320\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__33329\,
            I => \N__33317\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__33326\,
            I => \N__33314\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__33323\,
            I => \N__33311\
        );

    \I__6491\ : Span4Mux_v
    port map (
            O => \N__33320\,
            I => \N__33308\
        );

    \I__6490\ : Span4Mux_v
    port map (
            O => \N__33317\,
            I => \N__33305\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__33314\,
            I => \N__33302\
        );

    \I__6488\ : Odrv12
    port map (
            O => \N__33311\,
            I => \delay_measurement_inst.delay_tr_timer.N_435_i\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__33308\,
            I => \delay_measurement_inst.delay_tr_timer.N_435_i\
        );

    \I__6486\ : Odrv4
    port map (
            O => \N__33305\,
            I => \delay_measurement_inst.delay_tr_timer.N_435_i\
        );

    \I__6485\ : Odrv4
    port map (
            O => \N__33302\,
            I => \delay_measurement_inst.delay_tr_timer.N_435_i\
        );

    \I__6484\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33290\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__33290\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__6482\ : CascadeMux
    port map (
            O => \N__33287\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__33284\,
            I => \phase_controller_inst2.stoper_tr.running_1_sqmuxa_cascade_\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33274\
        );

    \I__6479\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33274\
        );

    \I__6478\ : InMux
    port map (
            O => \N__33279\,
            I => \N__33271\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__33274\,
            I => \N__33268\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__33271\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__6475\ : Odrv12
    port map (
            O => \N__33268\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__6474\ : InMux
    port map (
            O => \N__33263\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33253\
        );

    \I__6472\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33253\
        );

    \I__6471\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33250\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__33253\,
            I => \N__33247\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__33250\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__6468\ : Odrv12
    port map (
            O => \N__33247\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33242\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__6466\ : CascadeMux
    port map (
            O => \N__33239\,
            I => \N__33235\
        );

    \I__6465\ : CascadeMux
    port map (
            O => \N__33238\,
            I => \N__33232\
        );

    \I__6464\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33226\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33226\
        );

    \I__6462\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33223\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__33226\,
            I => \N__33220\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__33223\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__6459\ : Odrv12
    port map (
            O => \N__33220\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__6458\ : InMux
    port map (
            O => \N__33215\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__33212\,
            I => \N__33208\
        );

    \I__6456\ : CascadeMux
    port map (
            O => \N__33211\,
            I => \N__33205\
        );

    \I__6455\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33199\
        );

    \I__6454\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33199\
        );

    \I__6453\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33196\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__33199\,
            I => \N__33193\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__33196\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__6450\ : Odrv12
    port map (
            O => \N__33193\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__6449\ : InMux
    port map (
            O => \N__33188\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__6448\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33179\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33179\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__33179\,
            I => \N__33175\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33178\,
            I => \N__33172\
        );

    \I__6444\ : Span4Mux_v
    port map (
            O => \N__33175\,
            I => \N__33169\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__33172\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__6442\ : Odrv4
    port map (
            O => \N__33169\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33164\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__6440\ : CascadeMux
    port map (
            O => \N__33161\,
            I => \N__33158\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33158\,
            I => \N__33154\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33157\,
            I => \N__33151\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33154\,
            I => \N__33145\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__33151\,
            I => \N__33145\
        );

    \I__6435\ : InMux
    port map (
            O => \N__33150\,
            I => \N__33142\
        );

    \I__6434\ : Span4Mux_v
    port map (
            O => \N__33145\,
            I => \N__33139\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__33142\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__6432\ : Odrv4
    port map (
            O => \N__33139\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__6431\ : InMux
    port map (
            O => \N__33134\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__6430\ : CascadeMux
    port map (
            O => \N__33131\,
            I => \N__33127\
        );

    \I__6429\ : CascadeMux
    port map (
            O => \N__33130\,
            I => \N__33124\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33121\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33124\,
            I => \N__33118\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__33121\,
            I => \N__33112\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__33118\,
            I => \N__33112\
        );

    \I__6424\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33109\
        );

    \I__6423\ : Span4Mux_v
    port map (
            O => \N__33112\,
            I => \N__33106\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__33109\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__6421\ : Odrv4
    port map (
            O => \N__33106\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__6420\ : InMux
    port map (
            O => \N__33101\,
            I => \bfn_13_12_0_\
        );

    \I__6419\ : CascadeMux
    port map (
            O => \N__33098\,
            I => \N__33095\
        );

    \I__6418\ : InMux
    port map (
            O => \N__33095\,
            I => \N__33090\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33094\,
            I => \N__33087\
        );

    \I__6416\ : InMux
    port map (
            O => \N__33093\,
            I => \N__33084\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__33090\,
            I => \N__33079\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__33087\,
            I => \N__33079\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__33084\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__6412\ : Odrv12
    port map (
            O => \N__33079\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__6411\ : InMux
    port map (
            O => \N__33074\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__6410\ : InMux
    port map (
            O => \N__33071\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33062\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33062\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__33062\,
            I => \N__33058\
        );

    \I__6406\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33055\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__33058\,
            I => \N__33052\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__33055\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__33052\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__6402\ : InMux
    port map (
            O => \N__33047\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__6401\ : InMux
    port map (
            O => \N__33044\,
            I => \N__33038\
        );

    \I__6400\ : InMux
    port map (
            O => \N__33043\,
            I => \N__33038\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__33038\,
            I => \N__33034\
        );

    \I__6398\ : InMux
    port map (
            O => \N__33037\,
            I => \N__33031\
        );

    \I__6397\ : Span4Mux_v
    port map (
            O => \N__33034\,
            I => \N__33028\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__33031\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__33028\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33023\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__6393\ : CascadeMux
    port map (
            O => \N__33020\,
            I => \N__33016\
        );

    \I__6392\ : CascadeMux
    port map (
            O => \N__33019\,
            I => \N__33013\
        );

    \I__6391\ : InMux
    port map (
            O => \N__33016\,
            I => \N__33007\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33013\,
            I => \N__33007\
        );

    \I__6389\ : InMux
    port map (
            O => \N__33012\,
            I => \N__33004\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__33007\,
            I => \N__33001\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__33004\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__6386\ : Odrv12
    port map (
            O => \N__33001\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__6385\ : InMux
    port map (
            O => \N__32996\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__6384\ : CascadeMux
    port map (
            O => \N__32993\,
            I => \N__32989\
        );

    \I__6383\ : CascadeMux
    port map (
            O => \N__32992\,
            I => \N__32986\
        );

    \I__6382\ : InMux
    port map (
            O => \N__32989\,
            I => \N__32980\
        );

    \I__6381\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32980\
        );

    \I__6380\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32977\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__32980\,
            I => \N__32974\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__32977\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__6377\ : Odrv12
    port map (
            O => \N__32974\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__6376\ : InMux
    port map (
            O => \N__32969\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__6375\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32960\
        );

    \I__6374\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32960\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__32960\,
            I => \N__32956\
        );

    \I__6372\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32953\
        );

    \I__6371\ : Span4Mux_v
    port map (
            O => \N__32956\,
            I => \N__32950\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__32953\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__6369\ : Odrv4
    port map (
            O => \N__32950\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__6368\ : InMux
    port map (
            O => \N__32945\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__32942\,
            I => \N__32939\
        );

    \I__6366\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32935\
        );

    \I__6365\ : InMux
    port map (
            O => \N__32938\,
            I => \N__32932\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__32935\,
            I => \N__32926\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32926\
        );

    \I__6362\ : InMux
    port map (
            O => \N__32931\,
            I => \N__32923\
        );

    \I__6361\ : Span4Mux_v
    port map (
            O => \N__32926\,
            I => \N__32920\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__32923\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__32920\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__6358\ : InMux
    port map (
            O => \N__32915\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__6357\ : CascadeMux
    port map (
            O => \N__32912\,
            I => \N__32909\
        );

    \I__6356\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32905\
        );

    \I__6355\ : CascadeMux
    port map (
            O => \N__32908\,
            I => \N__32902\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__32905\,
            I => \N__32898\
        );

    \I__6353\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32895\
        );

    \I__6352\ : InMux
    port map (
            O => \N__32901\,
            I => \N__32892\
        );

    \I__6351\ : Sp12to4
    port map (
            O => \N__32898\,
            I => \N__32887\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__32895\,
            I => \N__32887\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__32892\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6348\ : Odrv12
    port map (
            O => \N__32887\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6347\ : InMux
    port map (
            O => \N__32882\,
            I => \bfn_13_11_0_\
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__32879\,
            I => \N__32876\
        );

    \I__6345\ : InMux
    port map (
            O => \N__32876\,
            I => \N__32873\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__32873\,
            I => \N__32868\
        );

    \I__6343\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32865\
        );

    \I__6342\ : InMux
    port map (
            O => \N__32871\,
            I => \N__32862\
        );

    \I__6341\ : Sp12to4
    port map (
            O => \N__32868\,
            I => \N__32857\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32857\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__32862\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6338\ : Odrv12
    port map (
            O => \N__32857\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6337\ : InMux
    port map (
            O => \N__32852\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__6336\ : InMux
    port map (
            O => \N__32849\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__6335\ : CascadeMux
    port map (
            O => \N__32846\,
            I => \N__32842\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32839\
        );

    \I__6333\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32836\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__32839\,
            I => \N__32830\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__32836\,
            I => \N__32830\
        );

    \I__6330\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32827\
        );

    \I__6329\ : Span4Mux_v
    port map (
            O => \N__32830\,
            I => \N__32824\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__32827\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__6327\ : Odrv4
    port map (
            O => \N__32824\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__6326\ : InMux
    port map (
            O => \N__32819\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__6325\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32810\
        );

    \I__6324\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32810\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__32810\,
            I => \N__32806\
        );

    \I__6322\ : InMux
    port map (
            O => \N__32809\,
            I => \N__32803\
        );

    \I__6321\ : Span4Mux_v
    port map (
            O => \N__32806\,
            I => \N__32800\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__32803\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__6319\ : Odrv4
    port map (
            O => \N__32800\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__6318\ : InMux
    port map (
            O => \N__32795\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__6317\ : CascadeMux
    port map (
            O => \N__32792\,
            I => \N__32788\
        );

    \I__6316\ : CascadeMux
    port map (
            O => \N__32791\,
            I => \N__32785\
        );

    \I__6315\ : InMux
    port map (
            O => \N__32788\,
            I => \N__32779\
        );

    \I__6314\ : InMux
    port map (
            O => \N__32785\,
            I => \N__32779\
        );

    \I__6313\ : InMux
    port map (
            O => \N__32784\,
            I => \N__32776\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__32779\,
            I => \N__32773\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__32776\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__6310\ : Odrv12
    port map (
            O => \N__32773\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__6309\ : InMux
    port map (
            O => \N__32768\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__6308\ : CascadeMux
    port map (
            O => \N__32765\,
            I => \N__32761\
        );

    \I__6307\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32757\
        );

    \I__6306\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32754\
        );

    \I__6305\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32751\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__32757\,
            I => \N__32746\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__32754\,
            I => \N__32746\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__32751\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__6301\ : Odrv12
    port map (
            O => \N__32746\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__6300\ : InMux
    port map (
            O => \N__32741\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__6299\ : InMux
    port map (
            O => \N__32738\,
            I => \N__32732\
        );

    \I__6298\ : InMux
    port map (
            O => \N__32737\,
            I => \N__32732\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__32732\,
            I => \N__32728\
        );

    \I__6296\ : InMux
    port map (
            O => \N__32731\,
            I => \N__32725\
        );

    \I__6295\ : Span4Mux_v
    port map (
            O => \N__32728\,
            I => \N__32722\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__32725\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__6293\ : Odrv4
    port map (
            O => \N__32722\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__6292\ : InMux
    port map (
            O => \N__32717\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__6291\ : CascadeMux
    port map (
            O => \N__32714\,
            I => \N__32710\
        );

    \I__6290\ : CascadeMux
    port map (
            O => \N__32713\,
            I => \N__32707\
        );

    \I__6289\ : InMux
    port map (
            O => \N__32710\,
            I => \N__32702\
        );

    \I__6288\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32702\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__32702\,
            I => \N__32698\
        );

    \I__6286\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32695\
        );

    \I__6285\ : Span4Mux_v
    port map (
            O => \N__32698\,
            I => \N__32692\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__32695\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__6283\ : Odrv4
    port map (
            O => \N__32692\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__6282\ : InMux
    port map (
            O => \N__32687\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__6281\ : CascadeMux
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__6280\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32677\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__32680\,
            I => \N__32674\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__32677\,
            I => \N__32670\
        );

    \I__6277\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32667\
        );

    \I__6276\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32664\
        );

    \I__6275\ : Sp12to4
    port map (
            O => \N__32670\,
            I => \N__32659\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__32667\,
            I => \N__32659\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__32664\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6272\ : Odrv12
    port map (
            O => \N__32659\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6271\ : InMux
    port map (
            O => \N__32654\,
            I => \bfn_13_10_0_\
        );

    \I__6270\ : CascadeMux
    port map (
            O => \N__32651\,
            I => \N__32648\
        );

    \I__6269\ : InMux
    port map (
            O => \N__32648\,
            I => \N__32645\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__32645\,
            I => \N__32640\
        );

    \I__6267\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32637\
        );

    \I__6266\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32634\
        );

    \I__6265\ : Sp12to4
    port map (
            O => \N__32640\,
            I => \N__32629\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__32637\,
            I => \N__32629\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__32634\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6262\ : Odrv12
    port map (
            O => \N__32629\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6261\ : InMux
    port map (
            O => \N__32624\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__6260\ : InMux
    port map (
            O => \N__32621\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__6259\ : InMux
    port map (
            O => \N__32618\,
            I => \bfn_13_8_0_\
        );

    \I__6258\ : InMux
    port map (
            O => \N__32615\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__6257\ : InMux
    port map (
            O => \N__32612\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__6256\ : InMux
    port map (
            O => \N__32609\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__6255\ : InMux
    port map (
            O => \N__32606\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__6254\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32579\
        );

    \I__6253\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32579\
        );

    \I__6252\ : InMux
    port map (
            O => \N__32601\,
            I => \N__32579\
        );

    \I__6251\ : InMux
    port map (
            O => \N__32600\,
            I => \N__32579\
        );

    \I__6250\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32570\
        );

    \I__6249\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32570\
        );

    \I__6248\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32570\
        );

    \I__6247\ : InMux
    port map (
            O => \N__32596\,
            I => \N__32570\
        );

    \I__6246\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32547\
        );

    \I__6245\ : InMux
    port map (
            O => \N__32594\,
            I => \N__32547\
        );

    \I__6244\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32547\
        );

    \I__6243\ : InMux
    port map (
            O => \N__32592\,
            I => \N__32547\
        );

    \I__6242\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32538\
        );

    \I__6241\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32538\
        );

    \I__6240\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32538\
        );

    \I__6239\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32538\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__32579\,
            I => \N__32535\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__32570\,
            I => \N__32532\
        );

    \I__6236\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32527\
        );

    \I__6235\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32527\
        );

    \I__6234\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32518\
        );

    \I__6233\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32518\
        );

    \I__6232\ : InMux
    port map (
            O => \N__32565\,
            I => \N__32518\
        );

    \I__6231\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32518\
        );

    \I__6230\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32509\
        );

    \I__6229\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32509\
        );

    \I__6228\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32509\
        );

    \I__6227\ : InMux
    port map (
            O => \N__32560\,
            I => \N__32509\
        );

    \I__6226\ : InMux
    port map (
            O => \N__32559\,
            I => \N__32500\
        );

    \I__6225\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32500\
        );

    \I__6224\ : InMux
    port map (
            O => \N__32557\,
            I => \N__32500\
        );

    \I__6223\ : InMux
    port map (
            O => \N__32556\,
            I => \N__32500\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__32547\,
            I => \N__32495\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__32538\,
            I => \N__32495\
        );

    \I__6220\ : Span4Mux_h
    port map (
            O => \N__32535\,
            I => \N__32490\
        );

    \I__6219\ : Span4Mux_h
    port map (
            O => \N__32532\,
            I => \N__32490\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__32527\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__32518\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__32509\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__32500\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__32495\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6213\ : Odrv4
    port map (
            O => \N__32490\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6212\ : InMux
    port map (
            O => \N__32477\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__6211\ : InMux
    port map (
            O => \N__32474\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__6210\ : InMux
    port map (
            O => \N__32471\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32468\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__6208\ : InMux
    port map (
            O => \N__32465\,
            I => \bfn_13_7_0_\
        );

    \I__6207\ : InMux
    port map (
            O => \N__32462\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32459\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__6205\ : InMux
    port map (
            O => \N__32456\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__6204\ : InMux
    port map (
            O => \N__32453\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__6203\ : InMux
    port map (
            O => \N__32450\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__6202\ : InMux
    port map (
            O => \N__32447\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__6201\ : InMux
    port map (
            O => \N__32444\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__6200\ : InMux
    port map (
            O => \N__32441\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__6199\ : InMux
    port map (
            O => \N__32438\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__6198\ : InMux
    port map (
            O => \N__32435\,
            I => \bfn_13_6_0_\
        );

    \I__6197\ : InMux
    port map (
            O => \N__32432\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__6196\ : InMux
    port map (
            O => \N__32429\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__6195\ : InMux
    port map (
            O => \N__32426\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__6194\ : InMux
    port map (
            O => \N__32423\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__6193\ : InMux
    port map (
            O => \N__32420\,
            I => \N__32415\
        );

    \I__6192\ : InMux
    port map (
            O => \N__32419\,
            I => \N__32412\
        );

    \I__6191\ : InMux
    port map (
            O => \N__32418\,
            I => \N__32409\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__32415\,
            I => \N__32403\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__32412\,
            I => \N__32403\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__32409\,
            I => \N__32400\
        );

    \I__6187\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32395\
        );

    \I__6186\ : Span4Mux_h
    port map (
            O => \N__32403\,
            I => \N__32392\
        );

    \I__6185\ : Span12Mux_h
    port map (
            O => \N__32400\,
            I => \N__32389\
        );

    \I__6184\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32386\
        );

    \I__6183\ : InMux
    port map (
            O => \N__32398\,
            I => \N__32383\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__32395\,
            I => \N__32378\
        );

    \I__6181\ : Span4Mux_h
    port map (
            O => \N__32392\,
            I => \N__32378\
        );

    \I__6180\ : Odrv12
    port map (
            O => \N__32389\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__32386\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__32383\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__6177\ : Odrv4
    port map (
            O => \N__32378\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__6176\ : InMux
    port map (
            O => \N__32369\,
            I => \N__32363\
        );

    \I__6175\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32363\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__32363\,
            I => \N__32358\
        );

    \I__6173\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32353\
        );

    \I__6172\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32353\
        );

    \I__6171\ : Odrv4
    port map (
            O => \N__32358\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__32353\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__6169\ : IoInMux
    port map (
            O => \N__32348\,
            I => \N__32345\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__32345\,
            I => \N__32342\
        );

    \I__6167\ : Span4Mux_s3_v
    port map (
            O => \N__32342\,
            I => \N__32339\
        );

    \I__6166\ : Span4Mux_v
    port map (
            O => \N__32339\,
            I => \N__32336\
        );

    \I__6165\ : Span4Mux_v
    port map (
            O => \N__32336\,
            I => \N__32332\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32329\
        );

    \I__6163\ : Odrv4
    port map (
            O => \N__32332\,
            I => \T45_c\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__32329\,
            I => \T45_c\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32321\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__32321\,
            I => \N__32318\
        );

    \I__6159\ : Span12Mux_v
    port map (
            O => \N__32318\,
            I => \N__32315\
        );

    \I__6158\ : Odrv12
    port map (
            O => \N__32315\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__6157\ : CEMux
    port map (
            O => \N__32312\,
            I => \N__32308\
        );

    \I__6156\ : CEMux
    port map (
            O => \N__32311\,
            I => \N__32304\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__32308\,
            I => \N__32301\
        );

    \I__6154\ : CEMux
    port map (
            O => \N__32307\,
            I => \N__32298\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__32304\,
            I => \N__32295\
        );

    \I__6152\ : Span4Mux_h
    port map (
            O => \N__32301\,
            I => \N__32289\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__32298\,
            I => \N__32289\
        );

    \I__6150\ : Span4Mux_v
    port map (
            O => \N__32295\,
            I => \N__32286\
        );

    \I__6149\ : CEMux
    port map (
            O => \N__32294\,
            I => \N__32283\
        );

    \I__6148\ : Odrv4
    port map (
            O => \N__32289\,
            I => \delay_measurement_inst.delay_hc_timer.N_433_i\
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__32286\,
            I => \delay_measurement_inst.delay_hc_timer.N_433_i\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__32283\,
            I => \delay_measurement_inst.delay_hc_timer.N_433_i\
        );

    \I__6145\ : InMux
    port map (
            O => \N__32276\,
            I => \N__32272\
        );

    \I__6144\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32269\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__32272\,
            I => \N__32262\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__32269\,
            I => \N__32262\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32268\,
            I => \N__32259\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32256\
        );

    \I__6139\ : Span12Mux_v
    port map (
            O => \N__32262\,
            I => \N__32253\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__32259\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__32256\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__6136\ : Odrv12
    port map (
            O => \N__32253\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32246\,
            I => \N__32241\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32238\
        );

    \I__6133\ : InMux
    port map (
            O => \N__32244\,
            I => \N__32235\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32241\,
            I => \N__32232\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__32238\,
            I => \N__32225\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__32235\,
            I => \N__32225\
        );

    \I__6129\ : Sp12to4
    port map (
            O => \N__32232\,
            I => \N__32225\
        );

    \I__6128\ : Span12Mux_v
    port map (
            O => \N__32225\,
            I => \N__32222\
        );

    \I__6127\ : Odrv12
    port map (
            O => \N__32222\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32219\,
            I => \N__32213\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32218\,
            I => \N__32210\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32217\,
            I => \N__32207\
        );

    \I__6123\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32204\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__32213\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__32210\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__32207\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__32204\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6118\ : InMux
    port map (
            O => \N__32195\,
            I => \bfn_13_5_0_\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32192\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32189\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__6115\ : InMux
    port map (
            O => \N__32186\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__6114\ : IoInMux
    port map (
            O => \N__32183\,
            I => \N__32180\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32180\,
            I => \N__32177\
        );

    \I__6112\ : IoSpan4Mux
    port map (
            O => \N__32177\,
            I => \N__32174\
        );

    \I__6111\ : Span4Mux_s1_v
    port map (
            O => \N__32174\,
            I => \N__32171\
        );

    \I__6110\ : Sp12to4
    port map (
            O => \N__32171\,
            I => \N__32168\
        );

    \I__6109\ : Span12Mux_v
    port map (
            O => \N__32168\,
            I => \N__32164\
        );

    \I__6108\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32161\
        );

    \I__6107\ : Odrv12
    port map (
            O => \N__32164\,
            I => \T12_c\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__32161\,
            I => \T12_c\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32153\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__32153\,
            I => \N__32150\
        );

    \I__6103\ : Span4Mux_v
    port map (
            O => \N__32150\,
            I => \N__32145\
        );

    \I__6102\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32140\
        );

    \I__6101\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32140\
        );

    \I__6100\ : Sp12to4
    port map (
            O => \N__32145\,
            I => \N__32133\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__32140\,
            I => \N__32133\
        );

    \I__6098\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32128\
        );

    \I__6097\ : InMux
    port map (
            O => \N__32138\,
            I => \N__32128\
        );

    \I__6096\ : Odrv12
    port map (
            O => \N__32133\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__32128\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__32123\,
            I => \N__32120\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32117\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__32117\,
            I => \N__32114\
        );

    \I__6091\ : Span4Mux_h
    port map (
            O => \N__32114\,
            I => \N__32108\
        );

    \I__6090\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32105\
        );

    \I__6089\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32102\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32099\
        );

    \I__6087\ : Span4Mux_h
    port map (
            O => \N__32108\,
            I => \N__32096\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__32105\,
            I => \N__32091\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__32102\,
            I => \N__32091\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32099\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__6083\ : Odrv4
    port map (
            O => \N__32096\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__6082\ : Odrv4
    port map (
            O => \N__32091\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__6081\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32081\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__32081\,
            I => \N__32078\
        );

    \I__6079\ : Span4Mux_v
    port map (
            O => \N__32078\,
            I => \N__32075\
        );

    \I__6078\ : Span4Mux_v
    port map (
            O => \N__32075\,
            I => \N__32071\
        );

    \I__6077\ : CascadeMux
    port map (
            O => \N__32074\,
            I => \N__32068\
        );

    \I__6076\ : Sp12to4
    port map (
            O => \N__32071\,
            I => \N__32064\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32059\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32059\
        );

    \I__6073\ : Span12Mux_h
    port map (
            O => \N__32064\,
            I => \N__32054\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32059\,
            I => \N__32054\
        );

    \I__6071\ : Span12Mux_v
    port map (
            O => \N__32054\,
            I => \N__32051\
        );

    \I__6070\ : Odrv12
    port map (
            O => \N__32051\,
            I => \il_max_comp2_D2\
        );

    \I__6069\ : CascadeMux
    port map (
            O => \N__32048\,
            I => \phase_controller_inst2.time_passed_RNI9M3O_cascade_\
        );

    \I__6068\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32042\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__32042\,
            I => \phase_controller_inst2.time_passed_RNI9M3O\
        );

    \I__6066\ : IoInMux
    port map (
            O => \N__32039\,
            I => \N__32036\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__32036\,
            I => \N__32033\
        );

    \I__6064\ : Span4Mux_s3_v
    port map (
            O => \N__32033\,
            I => \N__32030\
        );

    \I__6063\ : Span4Mux_h
    port map (
            O => \N__32030\,
            I => \N__32027\
        );

    \I__6062\ : Span4Mux_v
    port map (
            O => \N__32027\,
            I => \N__32024\
        );

    \I__6061\ : Span4Mux_v
    port map (
            O => \N__32024\,
            I => \N__32020\
        );

    \I__6060\ : InMux
    port map (
            O => \N__32023\,
            I => \N__32017\
        );

    \I__6059\ : Odrv4
    port map (
            O => \N__32020\,
            I => \T23_c\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__32017\,
            I => \T23_c\
        );

    \I__6057\ : CascadeMux
    port map (
            O => \N__32012\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6_cascade_\
        );

    \I__6056\ : InMux
    port map (
            O => \N__32009\,
            I => \N__32006\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__32006\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5\
        );

    \I__6054\ : InMux
    port map (
            O => \N__32003\,
            I => \N__31998\
        );

    \I__6053\ : InMux
    port map (
            O => \N__32002\,
            I => \N__31993\
        );

    \I__6052\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31993\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__31998\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__31993\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\
        );

    \I__6049\ : CascadeMux
    port map (
            O => \N__31988\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_\
        );

    \I__6048\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31982\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31979\
        );

    \I__6046\ : Span4Mux_h
    port map (
            O => \N__31979\,
            I => \N__31976\
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__31976\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31\
        );

    \I__6044\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31968\
        );

    \I__6043\ : InMux
    port map (
            O => \N__31972\,
            I => \N__31963\
        );

    \I__6042\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31963\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__31968\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__31963\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__31958\,
            I => \N__31955\
        );

    \I__6038\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31952\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__31952\,
            I => \N__31947\
        );

    \I__6036\ : InMux
    port map (
            O => \N__31951\,
            I => \N__31944\
        );

    \I__6035\ : InMux
    port map (
            O => \N__31950\,
            I => \N__31941\
        );

    \I__6034\ : Odrv4
    port map (
            O => \N__31947\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__31944\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__31941\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__6031\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31930\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__31933\,
            I => \N__31927\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__31930\,
            I => \N__31923\
        );

    \I__6028\ : InMux
    port map (
            O => \N__31927\,
            I => \N__31920\
        );

    \I__6027\ : InMux
    port map (
            O => \N__31926\,
            I => \N__31917\
        );

    \I__6026\ : Span4Mux_v
    port map (
            O => \N__31923\,
            I => \N__31914\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__31920\,
            I => \N__31911\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__31917\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__6023\ : Odrv4
    port map (
            O => \N__31914\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__6022\ : Odrv4
    port map (
            O => \N__31911\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__6021\ : InMux
    port map (
            O => \N__31904\,
            I => \N__31901\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__31901\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\
        );

    \I__6019\ : InMux
    port map (
            O => \N__31898\,
            I => \N__31895\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__31895\,
            I => \N__31891\
        );

    \I__6017\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31888\
        );

    \I__6016\ : Span4Mux_h
    port map (
            O => \N__31891\,
            I => \N__31881\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__31888\,
            I => \N__31881\
        );

    \I__6014\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31876\
        );

    \I__6013\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31876\
        );

    \I__6012\ : Odrv4
    port map (
            O => \N__31881\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__31876\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__31871\,
            I => \N__31868\
        );

    \I__6009\ : InMux
    port map (
            O => \N__31868\,
            I => \N__31865\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__31865\,
            I => \N__31862\
        );

    \I__6007\ : Span4Mux_v
    port map (
            O => \N__31862\,
            I => \N__31857\
        );

    \I__6006\ : InMux
    port map (
            O => \N__31861\,
            I => \N__31852\
        );

    \I__6005\ : InMux
    port map (
            O => \N__31860\,
            I => \N__31852\
        );

    \I__6004\ : Odrv4
    port map (
            O => \N__31857\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__31852\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\
        );

    \I__6002\ : CascadeMux
    port map (
            O => \N__31847\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__31844\,
            I => \N__31841\
        );

    \I__6000\ : InMux
    port map (
            O => \N__31841\,
            I => \N__31838\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__31838\,
            I => \N__31834\
        );

    \I__5998\ : InMux
    port map (
            O => \N__31837\,
            I => \N__31830\
        );

    \I__5997\ : Span4Mux_h
    port map (
            O => \N__31834\,
            I => \N__31827\
        );

    \I__5996\ : InMux
    port map (
            O => \N__31833\,
            I => \N__31824\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31830\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__31827\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__31824\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\
        );

    \I__5992\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31814\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__31814\,
            I => \N__31809\
        );

    \I__5990\ : InMux
    port map (
            O => \N__31813\,
            I => \N__31806\
        );

    \I__5989\ : InMux
    port map (
            O => \N__31812\,
            I => \N__31803\
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__31809\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__31806\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__31803\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__31796\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_\
        );

    \I__5984\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31788\
        );

    \I__5983\ : CascadeMux
    port map (
            O => \N__31792\,
            I => \N__31783\
        );

    \I__5982\ : InMux
    port map (
            O => \N__31791\,
            I => \N__31780\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__31788\,
            I => \N__31777\
        );

    \I__5980\ : InMux
    port map (
            O => \N__31787\,
            I => \N__31772\
        );

    \I__5979\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31772\
        );

    \I__5978\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31768\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__31780\,
            I => \N__31765\
        );

    \I__5976\ : Span4Mux_h
    port map (
            O => \N__31777\,
            I => \N__31762\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__31772\,
            I => \N__31759\
        );

    \I__5974\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31756\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__31768\,
            I => \N__31753\
        );

    \I__5972\ : Span4Mux_h
    port map (
            O => \N__31765\,
            I => \N__31750\
        );

    \I__5971\ : Span4Mux_v
    port map (
            O => \N__31762\,
            I => \N__31747\
        );

    \I__5970\ : Span4Mux_h
    port map (
            O => \N__31759\,
            I => \N__31740\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__31756\,
            I => \N__31740\
        );

    \I__5968\ : Span4Mux_h
    port map (
            O => \N__31753\,
            I => \N__31740\
        );

    \I__5967\ : Odrv4
    port map (
            O => \N__31750\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__5966\ : Odrv4
    port map (
            O => \N__31747\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__5965\ : Odrv4
    port map (
            O => \N__31740\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__5964\ : InMux
    port map (
            O => \N__31733\,
            I => \N__31729\
        );

    \I__5963\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31726\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__31729\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__31726\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__31721\,
            I => \N__31718\
        );

    \I__5959\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31715\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__31715\,
            I => \N__31711\
        );

    \I__5957\ : InMux
    port map (
            O => \N__31714\,
            I => \N__31708\
        );

    \I__5956\ : Odrv4
    port map (
            O => \N__31711\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__31708\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__5954\ : CascadeMux
    port map (
            O => \N__31703\,
            I => \N__31700\
        );

    \I__5953\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31697\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__31697\,
            I => \N__31694\
        );

    \I__5951\ : Span4Mux_v
    port map (
            O => \N__31694\,
            I => \N__31690\
        );

    \I__5950\ : InMux
    port map (
            O => \N__31693\,
            I => \N__31687\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__31690\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__31687\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__5947\ : InMux
    port map (
            O => \N__31682\,
            I => \N__31676\
        );

    \I__5946\ : InMux
    port map (
            O => \N__31681\,
            I => \N__31676\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__31676\,
            I => \N__31672\
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__31675\,
            I => \N__31669\
        );

    \I__5943\ : Span4Mux_v
    port map (
            O => \N__31672\,
            I => \N__31666\
        );

    \I__5942\ : InMux
    port map (
            O => \N__31669\,
            I => \N__31663\
        );

    \I__5941\ : Odrv4
    port map (
            O => \N__31666\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__31663\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\
        );

    \I__5939\ : IoInMux
    port map (
            O => \N__31658\,
            I => \N__31655\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31652\
        );

    \I__5937\ : Span4Mux_s2_v
    port map (
            O => \N__31652\,
            I => \N__31649\
        );

    \I__5936\ : Sp12to4
    port map (
            O => \N__31649\,
            I => \N__31646\
        );

    \I__5935\ : Span12Mux_h
    port map (
            O => \N__31646\,
            I => \N__31643\
        );

    \I__5934\ : Span12Mux_v
    port map (
            O => \N__31643\,
            I => \N__31639\
        );

    \I__5933\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31636\
        );

    \I__5932\ : Odrv12
    port map (
            O => \N__31639\,
            I => \T01_c\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__31636\,
            I => \T01_c\
        );

    \I__5930\ : CascadeMux
    port map (
            O => \N__31631\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15_cascade_\
        );

    \I__5929\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31625\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__31625\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__31622\,
            I => \N__31619\
        );

    \I__5926\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31616\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__31616\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31\
        );

    \I__5924\ : CascadeMux
    port map (
            O => \N__31613\,
            I => \N__31610\
        );

    \I__5923\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31607\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__31607\,
            I => \N__31604\
        );

    \I__5921\ : Span4Mux_h
    port map (
            O => \N__31604\,
            I => \N__31600\
        );

    \I__5920\ : InMux
    port map (
            O => \N__31603\,
            I => \N__31597\
        );

    \I__5919\ : Odrv4
    port map (
            O => \N__31600\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__31597\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__5917\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31588\
        );

    \I__5916\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31585\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__31588\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__31585\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__5913\ : InMux
    port map (
            O => \N__31580\,
            I => \N__31577\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__31577\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\
        );

    \I__5911\ : CascadeMux
    port map (
            O => \N__31574\,
            I => \N__31570\
        );

    \I__5910\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31567\
        );

    \I__5909\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31564\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__31567\,
            I => \N__31561\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__31564\,
            I => \N__31558\
        );

    \I__5906\ : Span4Mux_v
    port map (
            O => \N__31561\,
            I => \N__31555\
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__31558\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__31555\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__5903\ : CascadeMux
    port map (
            O => \N__31550\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4_cascade_\
        );

    \I__5902\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31544\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__31544\,
            I => \N__31541\
        );

    \I__5900\ : Span4Mux_v
    port map (
            O => \N__31541\,
            I => \N__31536\
        );

    \I__5899\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31531\
        );

    \I__5898\ : InMux
    port map (
            O => \N__31539\,
            I => \N__31531\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__31536\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__31531\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__5895\ : InMux
    port map (
            O => \N__31526\,
            I => \N__31523\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__31523\,
            I => \N__31520\
        );

    \I__5893\ : Span4Mux_h
    port map (
            O => \N__31520\,
            I => \N__31516\
        );

    \I__5892\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31513\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__31516\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__31513\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__31508\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1_cascade_\
        );

    \I__5888\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31502\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__31502\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__31499\,
            I => \N__31496\
        );

    \I__5885\ : InMux
    port map (
            O => \N__31496\,
            I => \N__31492\
        );

    \I__5884\ : InMux
    port map (
            O => \N__31495\,
            I => \N__31489\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__31492\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__31489\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__5881\ : InMux
    port map (
            O => \N__31484\,
            I => \N__31481\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__31481\,
            I => \N__31477\
        );

    \I__5879\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31474\
        );

    \I__5878\ : Odrv4
    port map (
            O => \N__31477\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__31474\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__31469\,
            I => \N__31466\
        );

    \I__5875\ : InMux
    port map (
            O => \N__31466\,
            I => \N__31463\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__31463\,
            I => \N__31459\
        );

    \I__5873\ : CascadeMux
    port map (
            O => \N__31462\,
            I => \N__31456\
        );

    \I__5872\ : Span4Mux_h
    port map (
            O => \N__31459\,
            I => \N__31453\
        );

    \I__5871\ : InMux
    port map (
            O => \N__31456\,
            I => \N__31450\
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__31453\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__31450\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__5868\ : CascadeMux
    port map (
            O => \N__31445\,
            I => \N__31442\
        );

    \I__5867\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31439\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__31439\,
            I => \N__31435\
        );

    \I__5865\ : InMux
    port map (
            O => \N__31438\,
            I => \N__31432\
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__31435\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__31432\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__31427\,
            I => \N__31424\
        );

    \I__5861\ : InMux
    port map (
            O => \N__31424\,
            I => \N__31420\
        );

    \I__5860\ : InMux
    port map (
            O => \N__31423\,
            I => \N__31417\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__31420\,
            I => \N__31414\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__31417\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\
        );

    \I__5857\ : Odrv4
    port map (
            O => \N__31414\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\
        );

    \I__5856\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31406\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__31406\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\
        );

    \I__5854\ : InMux
    port map (
            O => \N__31403\,
            I => \N__31400\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__31400\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3\
        );

    \I__5852\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31394\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__31394\,
            I => \N__31391\
        );

    \I__5850\ : Odrv4
    port map (
            O => \N__31391\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__5849\ : InMux
    port map (
            O => \N__31388\,
            I => \N__31385\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__31385\,
            I => \N__31380\
        );

    \I__5847\ : CascadeMux
    port map (
            O => \N__31384\,
            I => \N__31377\
        );

    \I__5846\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31374\
        );

    \I__5845\ : Span4Mux_h
    port map (
            O => \N__31380\,
            I => \N__31371\
        );

    \I__5844\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31368\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__31374\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__5842\ : Odrv4
    port map (
            O => \N__31371\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__31368\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__5840\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31358\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__31358\,
            I => \N__31354\
        );

    \I__5838\ : InMux
    port map (
            O => \N__31357\,
            I => \N__31350\
        );

    \I__5837\ : Span4Mux_v
    port map (
            O => \N__31354\,
            I => \N__31347\
        );

    \I__5836\ : InMux
    port map (
            O => \N__31353\,
            I => \N__31344\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__31350\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__31347\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__31344\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__31337\,
            I => \N__31334\
        );

    \I__5831\ : InMux
    port map (
            O => \N__31334\,
            I => \N__31330\
        );

    \I__5830\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31326\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__31330\,
            I => \N__31323\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31329\,
            I => \N__31320\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__31326\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__5826\ : Odrv4
    port map (
            O => \N__31323\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__31320\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31310\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31310\,
            I => \N__31306\
        );

    \I__5822\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31302\
        );

    \I__5821\ : Span4Mux_h
    port map (
            O => \N__31306\,
            I => \N__31299\
        );

    \I__5820\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31296\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__31302\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__5818\ : Odrv4
    port map (
            O => \N__31299\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__31296\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__5816\ : InMux
    port map (
            O => \N__31289\,
            I => \N__31286\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__31286\,
            I => \N__31282\
        );

    \I__5814\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31278\
        );

    \I__5813\ : Span4Mux_h
    port map (
            O => \N__31282\,
            I => \N__31275\
        );

    \I__5812\ : InMux
    port map (
            O => \N__31281\,
            I => \N__31272\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__31278\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__31275\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__31272\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5808\ : InMux
    port map (
            O => \N__31265\,
            I => \N__31262\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__31262\,
            I => \N__31259\
        );

    \I__5806\ : Odrv4
    port map (
            O => \N__31259\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__31256\,
            I => \N__31253\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31250\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__31250\,
            I => \N__31247\
        );

    \I__5802\ : Span4Mux_h
    port map (
            O => \N__31247\,
            I => \N__31242\
        );

    \I__5801\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31239\
        );

    \I__5800\ : InMux
    port map (
            O => \N__31245\,
            I => \N__31236\
        );

    \I__5799\ : Span4Mux_h
    port map (
            O => \N__31242\,
            I => \N__31232\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__31239\,
            I => \N__31227\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__31236\,
            I => \N__31227\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31224\
        );

    \I__5795\ : Span4Mux_h
    port map (
            O => \N__31232\,
            I => \N__31221\
        );

    \I__5794\ : Span4Mux_v
    port map (
            O => \N__31227\,
            I => \N__31218\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31224\,
            I => \elapsed_time_ns_1_RNIO0MD11_0_11\
        );

    \I__5792\ : Odrv4
    port map (
            O => \N__31221\,
            I => \elapsed_time_ns_1_RNIO0MD11_0_11\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__31218\,
            I => \elapsed_time_ns_1_RNIO0MD11_0_11\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31211\,
            I => \N__31206\
        );

    \I__5789\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31203\
        );

    \I__5788\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31200\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__31206\,
            I => \N__31197\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31203\,
            I => \N__31192\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31192\
        );

    \I__5784\ : Odrv4
    port map (
            O => \N__31197\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__31192\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\
        );

    \I__5782\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31184\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__31184\,
            I => \N__31179\
        );

    \I__5780\ : InMux
    port map (
            O => \N__31183\,
            I => \N__31176\
        );

    \I__5779\ : InMux
    port map (
            O => \N__31182\,
            I => \N__31173\
        );

    \I__5778\ : Odrv4
    port map (
            O => \N__31179\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__31176\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__31173\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__5775\ : InMux
    port map (
            O => \N__31166\,
            I => \N__31163\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__31163\,
            I => \N__31158\
        );

    \I__5773\ : InMux
    port map (
            O => \N__31162\,
            I => \N__31155\
        );

    \I__5772\ : InMux
    port map (
            O => \N__31161\,
            I => \N__31152\
        );

    \I__5771\ : Odrv4
    port map (
            O => \N__31158\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__31155\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__31152\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__5768\ : InMux
    port map (
            O => \N__31145\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__5767\ : InMux
    port map (
            O => \N__31142\,
            I => \bfn_12_12_0_\
        );

    \I__5766\ : InMux
    port map (
            O => \N__31139\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__5765\ : InMux
    port map (
            O => \N__31136\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__5764\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31129\
        );

    \I__5763\ : CascadeMux
    port map (
            O => \N__31132\,
            I => \N__31126\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__31129\,
            I => \N__31123\
        );

    \I__5761\ : InMux
    port map (
            O => \N__31126\,
            I => \N__31120\
        );

    \I__5760\ : Span4Mux_v
    port map (
            O => \N__31123\,
            I => \N__31114\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__31120\,
            I => \N__31114\
        );

    \I__5758\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31111\
        );

    \I__5757\ : Span4Mux_h
    port map (
            O => \N__31114\,
            I => \N__31108\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__31111\,
            I => \N__31105\
        );

    \I__5755\ : Odrv4
    port map (
            O => \N__31108\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__31105\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5753\ : InMux
    port map (
            O => \N__31100\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__5752\ : InMux
    port map (
            O => \N__31097\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__5751\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31091\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__31091\,
            I => \N__31087\
        );

    \I__5749\ : InMux
    port map (
            O => \N__31090\,
            I => \N__31084\
        );

    \I__5748\ : Span4Mux_v
    port map (
            O => \N__31087\,
            I => \N__31079\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__31084\,
            I => \N__31079\
        );

    \I__5746\ : Span4Mux_h
    port map (
            O => \N__31079\,
            I => \N__31075\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31078\,
            I => \N__31072\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__31075\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__31072\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5742\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31064\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__31064\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\
        );

    \I__5740\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31058\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__31058\,
            I => \N__31054\
        );

    \I__5738\ : InMux
    port map (
            O => \N__31057\,
            I => \N__31051\
        );

    \I__5737\ : Span4Mux_v
    port map (
            O => \N__31054\,
            I => \N__31046\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__31051\,
            I => \N__31046\
        );

    \I__5735\ : Span4Mux_h
    port map (
            O => \N__31046\,
            I => \N__31042\
        );

    \I__5734\ : InMux
    port map (
            O => \N__31045\,
            I => \N__31039\
        );

    \I__5733\ : Odrv4
    port map (
            O => \N__31042\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__31039\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__5731\ : InMux
    port map (
            O => \N__31034\,
            I => \N__31031\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__31031\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\
        );

    \I__5729\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31025\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__31025\,
            I => \N__31021\
        );

    \I__5727\ : InMux
    port map (
            O => \N__31024\,
            I => \N__31018\
        );

    \I__5726\ : Span4Mux_v
    port map (
            O => \N__31021\,
            I => \N__31013\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__31018\,
            I => \N__31013\
        );

    \I__5724\ : Span4Mux_h
    port map (
            O => \N__31013\,
            I => \N__31009\
        );

    \I__5723\ : InMux
    port map (
            O => \N__31012\,
            I => \N__31006\
        );

    \I__5722\ : Odrv4
    port map (
            O => \N__31009\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__31006\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__5720\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30998\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__30998\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\
        );

    \I__5718\ : InMux
    port map (
            O => \N__30995\,
            I => \N__30992\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__30992\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\
        );

    \I__5716\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30986\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__30986\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__5714\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30980\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__30980\,
            I => \N__30976\
        );

    \I__5712\ : InMux
    port map (
            O => \N__30979\,
            I => \N__30973\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__30976\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__30973\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__5709\ : InMux
    port map (
            O => \N__30968\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__5708\ : InMux
    port map (
            O => \N__30965\,
            I => \N__30962\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__30962\,
            I => \N__30958\
        );

    \I__5706\ : InMux
    port map (
            O => \N__30961\,
            I => \N__30955\
        );

    \I__5705\ : Odrv4
    port map (
            O => \N__30958\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__30955\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__5703\ : InMux
    port map (
            O => \N__30950\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__5702\ : InMux
    port map (
            O => \N__30947\,
            I => \N__30944\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__30944\,
            I => \N__30941\
        );

    \I__5700\ : Span4Mux_v
    port map (
            O => \N__30941\,
            I => \N__30938\
        );

    \I__5699\ : Span4Mux_h
    port map (
            O => \N__30938\,
            I => \N__30934\
        );

    \I__5698\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30931\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__30934\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__30931\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__5695\ : InMux
    port map (
            O => \N__30926\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__5694\ : CascadeMux
    port map (
            O => \N__30923\,
            I => \N__30919\
        );

    \I__5693\ : InMux
    port map (
            O => \N__30922\,
            I => \N__30916\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30913\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30908\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__30913\,
            I => \N__30908\
        );

    \I__5689\ : Span4Mux_h
    port map (
            O => \N__30908\,
            I => \N__30904\
        );

    \I__5688\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30901\
        );

    \I__5687\ : Odrv4
    port map (
            O => \N__30904\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__30901\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__5685\ : InMux
    port map (
            O => \N__30896\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__5684\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30889\
        );

    \I__5683\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30886\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__30889\,
            I => \N__30880\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__30886\,
            I => \N__30880\
        );

    \I__5680\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30877\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__30880\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__30877\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__5677\ : InMux
    port map (
            O => \N__30872\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__5676\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30865\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__30868\,
            I => \N__30862\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__30865\,
            I => \N__30859\
        );

    \I__5673\ : InMux
    port map (
            O => \N__30862\,
            I => \N__30856\
        );

    \I__5672\ : Span4Mux_h
    port map (
            O => \N__30859\,
            I => \N__30853\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__30856\,
            I => \N__30850\
        );

    \I__5670\ : Span4Mux_h
    port map (
            O => \N__30853\,
            I => \N__30846\
        );

    \I__5669\ : Span4Mux_h
    port map (
            O => \N__30850\,
            I => \N__30843\
        );

    \I__5668\ : InMux
    port map (
            O => \N__30849\,
            I => \N__30840\
        );

    \I__5667\ : Odrv4
    port map (
            O => \N__30846\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__30843\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__30840\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__5664\ : InMux
    port map (
            O => \N__30833\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__30830\,
            I => \N__30826\
        );

    \I__5662\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30823\
        );

    \I__5661\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30820\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__30823\,
            I => \N__30815\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__30820\,
            I => \N__30815\
        );

    \I__5658\ : Span4Mux_h
    port map (
            O => \N__30815\,
            I => \N__30811\
        );

    \I__5657\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30808\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__30811\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__30808\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__30803\,
            I => \N__30800\
        );

    \I__5653\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30797\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__30797\,
            I => \N__30794\
        );

    \I__5651\ : Span12Mux_s8_h
    port map (
            O => \N__30794\,
            I => \N__30791\
        );

    \I__5650\ : Odrv12
    port map (
            O => \N__30791\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__5649\ : InMux
    port map (
            O => \N__30788\,
            I => \N__30785\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__30785\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__30782\,
            I => \N__30778\
        );

    \I__5646\ : CascadeMux
    port map (
            O => \N__30781\,
            I => \N__30775\
        );

    \I__5645\ : InMux
    port map (
            O => \N__30778\,
            I => \N__30772\
        );

    \I__5644\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30769\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__30772\,
            I => \N__30764\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__30769\,
            I => \N__30761\
        );

    \I__5641\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30758\
        );

    \I__5640\ : InMux
    port map (
            O => \N__30767\,
            I => \N__30755\
        );

    \I__5639\ : Span4Mux_v
    port map (
            O => \N__30764\,
            I => \N__30752\
        );

    \I__5638\ : Span4Mux_v
    port map (
            O => \N__30761\,
            I => \N__30747\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__30758\,
            I => \N__30747\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__30755\,
            I => \N__30741\
        );

    \I__5635\ : Span4Mux_h
    port map (
            O => \N__30752\,
            I => \N__30741\
        );

    \I__5634\ : Span4Mux_h
    port map (
            O => \N__30747\,
            I => \N__30738\
        );

    \I__5633\ : InMux
    port map (
            O => \N__30746\,
            I => \N__30735\
        );

    \I__5632\ : Odrv4
    port map (
            O => \N__30741\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__5631\ : Odrv4
    port map (
            O => \N__30738\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__30735\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__5629\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30725\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__30725\,
            I => \N__30722\
        );

    \I__5627\ : Span4Mux_v
    port map (
            O => \N__30722\,
            I => \N__30719\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__30719\,
            I => \current_shift_inst.PI_CTRL.integrator_i_8\
        );

    \I__5625\ : InMux
    port map (
            O => \N__30716\,
            I => \N__30713\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__30713\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\
        );

    \I__5623\ : InMux
    port map (
            O => \N__30710\,
            I => \N__30707\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__30707\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\
        );

    \I__5621\ : InMux
    port map (
            O => \N__30704\,
            I => \N__30701\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__30701\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\
        );

    \I__5619\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30693\
        );

    \I__5618\ : InMux
    port map (
            O => \N__30697\,
            I => \N__30690\
        );

    \I__5617\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30687\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__30693\,
            I => \N__30684\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__30690\,
            I => \N__30681\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__30687\,
            I => \N__30676\
        );

    \I__5613\ : Span4Mux_h
    port map (
            O => \N__30684\,
            I => \N__30671\
        );

    \I__5612\ : Span4Mux_h
    port map (
            O => \N__30681\,
            I => \N__30671\
        );

    \I__5611\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30668\
        );

    \I__5610\ : InMux
    port map (
            O => \N__30679\,
            I => \N__30665\
        );

    \I__5609\ : Span4Mux_v
    port map (
            O => \N__30676\,
            I => \N__30662\
        );

    \I__5608\ : Odrv4
    port map (
            O => \N__30671\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__30668\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__30665\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__30662\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5604\ : InMux
    port map (
            O => \N__30653\,
            I => \N__30650\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__30650\,
            I => \N__30647\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__30647\,
            I => \current_shift_inst.PI_CTRL.integrator_i_21\
        );

    \I__5601\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30641\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__30641\,
            I => \N__30636\
        );

    \I__5599\ : InMux
    port map (
            O => \N__30640\,
            I => \N__30633\
        );

    \I__5598\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30630\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__30636\,
            I => \N__30627\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__30633\,
            I => \N__30624\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__30630\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5594\ : Odrv4
    port map (
            O => \N__30627\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__30624\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5592\ : IoInMux
    port map (
            O => \N__30617\,
            I => \N__30614\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__30614\,
            I => \N__30611\
        );

    \I__5590\ : Span4Mux_s2_v
    port map (
            O => \N__30611\,
            I => \N__30608\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__30608\,
            I => \N__30605\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__30605\,
            I => \N__30602\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__30602\,
            I => \delay_measurement_inst.delay_hc_timer.N_432_i\
        );

    \I__5586\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30596\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__30596\,
            I => \N__30593\
        );

    \I__5584\ : Span4Mux_h
    port map (
            O => \N__30593\,
            I => \N__30590\
        );

    \I__5583\ : Odrv4
    port map (
            O => \N__30590\,
            I => il_min_comp1_c
        );

    \I__5582\ : InMux
    port map (
            O => \N__30587\,
            I => \N__30584\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__30584\,
            I => \il_min_comp1_D1\
        );

    \I__5580\ : ClkMux
    port map (
            O => \N__30581\,
            I => \N__30575\
        );

    \I__5579\ : ClkMux
    port map (
            O => \N__30580\,
            I => \N__30575\
        );

    \I__5578\ : GlobalMux
    port map (
            O => \N__30575\,
            I => \N__30572\
        );

    \I__5577\ : gio2CtrlBuf
    port map (
            O => \N__30572\,
            I => delay_hc_input_c_g
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__30569\,
            I => \N__30565\
        );

    \I__5575\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30562\
        );

    \I__5574\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30559\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__30562\,
            I => \N__30554\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30551\
        );

    \I__5571\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30548\
        );

    \I__5570\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30545\
        );

    \I__5569\ : Span4Mux_h
    port map (
            O => \N__30554\,
            I => \N__30542\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__30551\,
            I => \N__30539\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__30548\,
            I => \N__30534\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__30545\,
            I => \N__30534\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__30542\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__30539\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__5563\ : Odrv12
    port map (
            O => \N__30534\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__5562\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30524\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__30524\,
            I => \N__30521\
        );

    \I__5560\ : Odrv12
    port map (
            O => \N__30521\,
            I => \current_shift_inst.PI_CTRL.integrator_i_1\
        );

    \I__5559\ : CascadeMux
    port map (
            O => \N__30518\,
            I => \N__30515\
        );

    \I__5558\ : InMux
    port map (
            O => \N__30515\,
            I => \N__30511\
        );

    \I__5557\ : InMux
    port map (
            O => \N__30514\,
            I => \N__30508\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__30511\,
            I => \N__30503\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__30508\,
            I => \N__30503\
        );

    \I__5554\ : Odrv12
    port map (
            O => \N__30503\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_12\
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__30500\,
            I => \N__30496\
        );

    \I__5552\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30492\
        );

    \I__5551\ : InMux
    port map (
            O => \N__30496\,
            I => \N__30489\
        );

    \I__5550\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30486\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__30492\,
            I => \N__30483\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__30489\,
            I => \N__30480\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__30486\,
            I => \N__30477\
        );

    \I__5546\ : Span4Mux_h
    port map (
            O => \N__30483\,
            I => \N__30472\
        );

    \I__5545\ : Span4Mux_v
    port map (
            O => \N__30480\,
            I => \N__30469\
        );

    \I__5544\ : Span4Mux_v
    port map (
            O => \N__30477\,
            I => \N__30466\
        );

    \I__5543\ : InMux
    port map (
            O => \N__30476\,
            I => \N__30463\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30460\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__30472\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5540\ : Odrv4
    port map (
            O => \N__30469\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5539\ : Odrv4
    port map (
            O => \N__30466\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__30463\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__30460\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5536\ : InMux
    port map (
            O => \N__30449\,
            I => \N__30446\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__30446\,
            I => \N__30443\
        );

    \I__5534\ : Span4Mux_h
    port map (
            O => \N__30443\,
            I => \N__30440\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__30440\,
            I => \current_shift_inst.PI_CTRL.integrator_i_24\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__30437\,
            I => \N__30433\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__30436\,
            I => \N__30430\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30433\,
            I => \N__30424\
        );

    \I__5529\ : InMux
    port map (
            O => \N__30430\,
            I => \N__30424\
        );

    \I__5528\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30421\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30418\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__30421\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__5525\ : Odrv12
    port map (
            O => \N__30418\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__5524\ : InMux
    port map (
            O => \N__30413\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__30410\,
            I => \N__30406\
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__30409\,
            I => \N__30403\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30397\
        );

    \I__5520\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30397\
        );

    \I__5519\ : InMux
    port map (
            O => \N__30402\,
            I => \N__30394\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30391\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__30394\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__5516\ : Odrv12
    port map (
            O => \N__30391\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__5515\ : InMux
    port map (
            O => \N__30386\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__5514\ : CascadeMux
    port map (
            O => \N__30383\,
            I => \N__30380\
        );

    \I__5513\ : InMux
    port map (
            O => \N__30380\,
            I => \N__30375\
        );

    \I__5512\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30372\
        );

    \I__5511\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30369\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__30375\,
            I => \N__30364\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__30372\,
            I => \N__30364\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__30369\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__5507\ : Odrv12
    port map (
            O => \N__30364\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__5506\ : InMux
    port map (
            O => \N__30359\,
            I => \bfn_11_22_0_\
        );

    \I__5505\ : InMux
    port map (
            O => \N__30356\,
            I => \N__30352\
        );

    \I__5504\ : InMux
    port map (
            O => \N__30355\,
            I => \N__30349\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__30352\,
            I => \N__30343\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__30349\,
            I => \N__30343\
        );

    \I__5501\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30340\
        );

    \I__5500\ : Span4Mux_v
    port map (
            O => \N__30343\,
            I => \N__30337\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__30340\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__5498\ : Odrv4
    port map (
            O => \N__30337\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__5497\ : InMux
    port map (
            O => \N__30332\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__5496\ : CascadeMux
    port map (
            O => \N__30329\,
            I => \N__30326\
        );

    \I__5495\ : InMux
    port map (
            O => \N__30326\,
            I => \N__30322\
        );

    \I__5494\ : InMux
    port map (
            O => \N__30325\,
            I => \N__30319\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__30322\,
            I => \N__30313\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__30319\,
            I => \N__30313\
        );

    \I__5491\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30310\
        );

    \I__5490\ : Span4Mux_h
    port map (
            O => \N__30313\,
            I => \N__30307\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30310\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__30307\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__5487\ : InMux
    port map (
            O => \N__30302\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__5486\ : CascadeMux
    port map (
            O => \N__30299\,
            I => \N__30295\
        );

    \I__5485\ : CascadeMux
    port map (
            O => \N__30298\,
            I => \N__30292\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30286\
        );

    \I__5483\ : InMux
    port map (
            O => \N__30292\,
            I => \N__30286\
        );

    \I__5482\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30283\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__30286\,
            I => \N__30280\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30283\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__5479\ : Odrv12
    port map (
            O => \N__30280\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__5478\ : InMux
    port map (
            O => \N__30275\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30272\,
            I => \N__30268\
        );

    \I__5476\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30265\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30268\,
            I => \N__30262\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__30265\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__5473\ : Odrv12
    port map (
            O => \N__30262\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__5472\ : InMux
    port map (
            O => \N__30257\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__5471\ : InMux
    port map (
            O => \N__30254\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__5470\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30247\
        );

    \I__5469\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30244\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__30247\,
            I => \N__30241\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__30244\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__5466\ : Odrv12
    port map (
            O => \N__30241\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__5465\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30204\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30204\
        );

    \I__5463\ : InMux
    port map (
            O => \N__30234\,
            I => \N__30204\
        );

    \I__5462\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30204\
        );

    \I__5461\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30195\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30231\,
            I => \N__30195\
        );

    \I__5459\ : InMux
    port map (
            O => \N__30230\,
            I => \N__30195\
        );

    \I__5458\ : InMux
    port map (
            O => \N__30229\,
            I => \N__30195\
        );

    \I__5457\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30180\
        );

    \I__5456\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30180\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30226\,
            I => \N__30180\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30225\,
            I => \N__30180\
        );

    \I__5453\ : InMux
    port map (
            O => \N__30224\,
            I => \N__30171\
        );

    \I__5452\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30171\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30222\,
            I => \N__30171\
        );

    \I__5450\ : InMux
    port map (
            O => \N__30221\,
            I => \N__30171\
        );

    \I__5449\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30162\
        );

    \I__5448\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30162\
        );

    \I__5447\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30162\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30162\
        );

    \I__5445\ : InMux
    port map (
            O => \N__30216\,
            I => \N__30153\
        );

    \I__5444\ : InMux
    port map (
            O => \N__30215\,
            I => \N__30153\
        );

    \I__5443\ : InMux
    port map (
            O => \N__30214\,
            I => \N__30153\
        );

    \I__5442\ : InMux
    port map (
            O => \N__30213\,
            I => \N__30153\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__30204\,
            I => \N__30150\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__30195\,
            I => \N__30147\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30142\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30193\,
            I => \N__30142\
        );

    \I__5437\ : InMux
    port map (
            O => \N__30192\,
            I => \N__30133\
        );

    \I__5436\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30133\
        );

    \I__5435\ : InMux
    port map (
            O => \N__30190\,
            I => \N__30133\
        );

    \I__5434\ : InMux
    port map (
            O => \N__30189\,
            I => \N__30133\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__30180\,
            I => \N__30130\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__30171\,
            I => \N__30119\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30162\,
            I => \N__30119\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__30153\,
            I => \N__30119\
        );

    \I__5429\ : Span4Mux_h
    port map (
            O => \N__30150\,
            I => \N__30119\
        );

    \I__5428\ : Span4Mux_h
    port map (
            O => \N__30147\,
            I => \N__30119\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__30142\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__30133\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__30130\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5424\ : Odrv4
    port map (
            O => \N__30119\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__30110\,
            I => \N__30107\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30103\
        );

    \I__5421\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30100\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__30103\,
            I => \N__30094\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__30100\,
            I => \N__30094\
        );

    \I__5418\ : InMux
    port map (
            O => \N__30099\,
            I => \N__30091\
        );

    \I__5417\ : Span4Mux_v
    port map (
            O => \N__30094\,
            I => \N__30088\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__30091\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__5415\ : Odrv4
    port map (
            O => \N__30088\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__5414\ : InMux
    port map (
            O => \N__30083\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__5413\ : InMux
    port map (
            O => \N__30080\,
            I => \N__30074\
        );

    \I__5412\ : InMux
    port map (
            O => \N__30079\,
            I => \N__30074\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__30074\,
            I => \N__30070\
        );

    \I__5410\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30067\
        );

    \I__5409\ : Span4Mux_v
    port map (
            O => \N__30070\,
            I => \N__30064\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__30067\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__30064\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__5406\ : InMux
    port map (
            O => \N__30059\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__5405\ : CascadeMux
    port map (
            O => \N__30056\,
            I => \N__30053\
        );

    \I__5404\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30049\
        );

    \I__5403\ : InMux
    port map (
            O => \N__30052\,
            I => \N__30046\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__30049\,
            I => \N__30042\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__30046\,
            I => \N__30039\
        );

    \I__5400\ : InMux
    port map (
            O => \N__30045\,
            I => \N__30036\
        );

    \I__5399\ : Span4Mux_v
    port map (
            O => \N__30042\,
            I => \N__30031\
        );

    \I__5398\ : Span4Mux_v
    port map (
            O => \N__30039\,
            I => \N__30031\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__30036\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__5396\ : Odrv4
    port map (
            O => \N__30031\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30026\,
            I => \bfn_11_21_0_\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__30023\,
            I => \N__30019\
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__30022\,
            I => \N__30016\
        );

    \I__5392\ : InMux
    port map (
            O => \N__30019\,
            I => \N__30013\
        );

    \I__5391\ : InMux
    port map (
            O => \N__30016\,
            I => \N__30010\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__30013\,
            I => \N__30004\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__30010\,
            I => \N__30004\
        );

    \I__5388\ : InMux
    port map (
            O => \N__30009\,
            I => \N__30001\
        );

    \I__5387\ : Span4Mux_v
    port map (
            O => \N__30004\,
            I => \N__29998\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__30001\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__5385\ : Odrv4
    port map (
            O => \N__29998\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__5384\ : InMux
    port map (
            O => \N__29993\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__29990\,
            I => \N__29987\
        );

    \I__5382\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29983\
        );

    \I__5381\ : InMux
    port map (
            O => \N__29986\,
            I => \N__29980\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__29983\,
            I => \N__29974\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__29980\,
            I => \N__29974\
        );

    \I__5378\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29971\
        );

    \I__5377\ : Span4Mux_h
    port map (
            O => \N__29974\,
            I => \N__29968\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__29971\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__29968\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__5374\ : InMux
    port map (
            O => \N__29963\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__5373\ : InMux
    port map (
            O => \N__29960\,
            I => \N__29953\
        );

    \I__5372\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29953\
        );

    \I__5371\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29950\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__29953\,
            I => \N__29947\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__29950\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__5368\ : Odrv12
    port map (
            O => \N__29947\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__5367\ : InMux
    port map (
            O => \N__29942\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__5366\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29932\
        );

    \I__5365\ : InMux
    port map (
            O => \N__29938\,
            I => \N__29932\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29937\,
            I => \N__29929\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__29932\,
            I => \N__29926\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__29929\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__5361\ : Odrv12
    port map (
            O => \N__29926\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__5360\ : InMux
    port map (
            O => \N__29921\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__29918\,
            I => \N__29914\
        );

    \I__5358\ : InMux
    port map (
            O => \N__29917\,
            I => \N__29910\
        );

    \I__5357\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29907\
        );

    \I__5356\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29904\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__29910\,
            I => \N__29899\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__29907\,
            I => \N__29899\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__29904\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__5352\ : Odrv12
    port map (
            O => \N__29899\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__5351\ : InMux
    port map (
            O => \N__29894\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__5350\ : InMux
    port map (
            O => \N__29891\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__5349\ : CascadeMux
    port map (
            O => \N__29888\,
            I => \N__29885\
        );

    \I__5348\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29881\
        );

    \I__5347\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29878\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29872\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__29878\,
            I => \N__29872\
        );

    \I__5344\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29869\
        );

    \I__5343\ : Span4Mux_v
    port map (
            O => \N__29872\,
            I => \N__29866\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__29869\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__5341\ : Odrv4
    port map (
            O => \N__29866\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__5340\ : InMux
    port map (
            O => \N__29861\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__5339\ : InMux
    port map (
            O => \N__29858\,
            I => \N__29852\
        );

    \I__5338\ : InMux
    port map (
            O => \N__29857\,
            I => \N__29852\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__29852\,
            I => \N__29848\
        );

    \I__5336\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29845\
        );

    \I__5335\ : Span4Mux_v
    port map (
            O => \N__29848\,
            I => \N__29842\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__29845\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__29842\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__5332\ : InMux
    port map (
            O => \N__29837\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__5331\ : CascadeMux
    port map (
            O => \N__29834\,
            I => \N__29831\
        );

    \I__5330\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29828\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29823\
        );

    \I__5328\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29820\
        );

    \I__5327\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29817\
        );

    \I__5326\ : Span4Mux_v
    port map (
            O => \N__29823\,
            I => \N__29814\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29811\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__29817\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__29814\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__5322\ : Odrv12
    port map (
            O => \N__29811\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__5321\ : InMux
    port map (
            O => \N__29804\,
            I => \bfn_11_20_0_\
        );

    \I__5320\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29797\
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__29800\,
            I => \N__29794\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__29797\,
            I => \N__29790\
        );

    \I__5317\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29787\
        );

    \I__5316\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29784\
        );

    \I__5315\ : Span4Mux_h
    port map (
            O => \N__29790\,
            I => \N__29781\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__29787\,
            I => \N__29778\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__29784\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__29781\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__5311\ : Odrv12
    port map (
            O => \N__29778\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__5310\ : InMux
    port map (
            O => \N__29771\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__5309\ : InMux
    port map (
            O => \N__29768\,
            I => \N__29762\
        );

    \I__5308\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29762\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__29762\,
            I => \N__29758\
        );

    \I__5306\ : InMux
    port map (
            O => \N__29761\,
            I => \N__29755\
        );

    \I__5305\ : Span4Mux_v
    port map (
            O => \N__29758\,
            I => \N__29752\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__29755\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__5303\ : Odrv4
    port map (
            O => \N__29752\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__5302\ : InMux
    port map (
            O => \N__29747\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__5301\ : CascadeMux
    port map (
            O => \N__29744\,
            I => \N__29740\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__29743\,
            I => \N__29737\
        );

    \I__5299\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29731\
        );

    \I__5298\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29731\
        );

    \I__5297\ : InMux
    port map (
            O => \N__29736\,
            I => \N__29728\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__29731\,
            I => \N__29725\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__29728\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__5294\ : Odrv12
    port map (
            O => \N__29725\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__5293\ : InMux
    port map (
            O => \N__29720\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__5292\ : CascadeMux
    port map (
            O => \N__29717\,
            I => \N__29713\
        );

    \I__5291\ : CascadeMux
    port map (
            O => \N__29716\,
            I => \N__29710\
        );

    \I__5290\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29704\
        );

    \I__5289\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29704\
        );

    \I__5288\ : InMux
    port map (
            O => \N__29709\,
            I => \N__29701\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__29704\,
            I => \N__29698\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__29701\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__5285\ : Odrv12
    port map (
            O => \N__29698\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__5284\ : InMux
    port map (
            O => \N__29693\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__5283\ : CascadeMux
    port map (
            O => \N__29690\,
            I => \N__29687\
        );

    \I__5282\ : InMux
    port map (
            O => \N__29687\,
            I => \N__29683\
        );

    \I__5281\ : InMux
    port map (
            O => \N__29686\,
            I => \N__29680\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__29683\,
            I => \N__29674\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__29680\,
            I => \N__29674\
        );

    \I__5278\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29671\
        );

    \I__5277\ : Span4Mux_v
    port map (
            O => \N__29674\,
            I => \N__29668\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__29671\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__5275\ : Odrv4
    port map (
            O => \N__29668\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__5274\ : InMux
    port map (
            O => \N__29663\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__5273\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29657\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__29657\,
            I => \N__29654\
        );

    \I__5271\ : Span4Mux_h
    port map (
            O => \N__29654\,
            I => \N__29650\
        );

    \I__5270\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29647\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__29650\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__29647\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__5267\ : InMux
    port map (
            O => \N__29642\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__5266\ : InMux
    port map (
            O => \N__29639\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__5265\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29632\
        );

    \I__5264\ : InMux
    port map (
            O => \N__29635\,
            I => \N__29628\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__29632\,
            I => \N__29625\
        );

    \I__5262\ : InMux
    port map (
            O => \N__29631\,
            I => \N__29622\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__29628\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__5260\ : Odrv12
    port map (
            O => \N__29625\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__29622\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__5258\ : InMux
    port map (
            O => \N__29615\,
            I => \bfn_11_19_0_\
        );

    \I__5257\ : InMux
    port map (
            O => \N__29612\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__5256\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29605\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__29608\,
            I => \N__29602\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__29605\,
            I => \N__29598\
        );

    \I__5253\ : InMux
    port map (
            O => \N__29602\,
            I => \N__29595\
        );

    \I__5252\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29592\
        );

    \I__5251\ : Span4Mux_h
    port map (
            O => \N__29598\,
            I => \N__29589\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__29595\,
            I => \N__29586\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__29592\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__5248\ : Odrv4
    port map (
            O => \N__29589\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__5247\ : Odrv12
    port map (
            O => \N__29586\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__5246\ : InMux
    port map (
            O => \N__29579\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__29576\,
            I => \N__29572\
        );

    \I__5244\ : InMux
    port map (
            O => \N__29575\,
            I => \N__29569\
        );

    \I__5243\ : InMux
    port map (
            O => \N__29572\,
            I => \N__29566\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__29569\,
            I => \N__29560\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__29566\,
            I => \N__29560\
        );

    \I__5240\ : InMux
    port map (
            O => \N__29565\,
            I => \N__29557\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__29560\,
            I => \N__29554\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__29557\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__29554\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__5236\ : InMux
    port map (
            O => \N__29549\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__5235\ : CascadeMux
    port map (
            O => \N__29546\,
            I => \N__29542\
        );

    \I__5234\ : CascadeMux
    port map (
            O => \N__29545\,
            I => \N__29539\
        );

    \I__5233\ : InMux
    port map (
            O => \N__29542\,
            I => \N__29533\
        );

    \I__5232\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29533\
        );

    \I__5231\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29530\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__29533\,
            I => \N__29527\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__29530\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__5228\ : Odrv12
    port map (
            O => \N__29527\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__5227\ : InMux
    port map (
            O => \N__29522\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__29519\,
            I => \N__29515\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__29518\,
            I => \N__29512\
        );

    \I__5224\ : InMux
    port map (
            O => \N__29515\,
            I => \N__29507\
        );

    \I__5223\ : InMux
    port map (
            O => \N__29512\,
            I => \N__29507\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__29507\,
            I => \N__29503\
        );

    \I__5221\ : InMux
    port map (
            O => \N__29506\,
            I => \N__29500\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__29503\,
            I => \N__29497\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__29500\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__5218\ : Odrv4
    port map (
            O => \N__29497\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__5217\ : InMux
    port map (
            O => \N__29492\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__5216\ : InMux
    port map (
            O => \N__29489\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__5215\ : InMux
    port map (
            O => \N__29486\,
            I => \N__29483\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__29483\,
            I => \N__29479\
        );

    \I__5213\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29476\
        );

    \I__5212\ : Odrv4
    port map (
            O => \N__29479\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__29476\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__5210\ : InMux
    port map (
            O => \N__29471\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__5209\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29465\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__29465\,
            I => \N__29461\
        );

    \I__5207\ : InMux
    port map (
            O => \N__29464\,
            I => \N__29458\
        );

    \I__5206\ : Odrv4
    port map (
            O => \N__29461\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__29458\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5204\ : InMux
    port map (
            O => \N__29453\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__5203\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29447\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__29447\,
            I => \N__29443\
        );

    \I__5201\ : CascadeMux
    port map (
            O => \N__29446\,
            I => \N__29440\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__29443\,
            I => \N__29437\
        );

    \I__5199\ : InMux
    port map (
            O => \N__29440\,
            I => \N__29434\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__29437\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__29434\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29429\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__29426\,
            I => \N__29423\
        );

    \I__5194\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29420\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29417\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__29417\,
            I => \N__29413\
        );

    \I__5191\ : InMux
    port map (
            O => \N__29416\,
            I => \N__29410\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__29413\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__29410\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29405\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__5187\ : CascadeMux
    port map (
            O => \N__29402\,
            I => \N__29399\
        );

    \I__5186\ : InMux
    port map (
            O => \N__29399\,
            I => \N__29396\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__29396\,
            I => \N__29393\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__29393\,
            I => \N__29390\
        );

    \I__5183\ : Span4Mux_v
    port map (
            O => \N__29390\,
            I => \N__29386\
        );

    \I__5182\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29383\
        );

    \I__5181\ : Odrv4
    port map (
            O => \N__29386\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__29383\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29378\,
            I => \bfn_11_18_0_\
        );

    \I__5178\ : CascadeMux
    port map (
            O => \N__29375\,
            I => \N__29372\
        );

    \I__5177\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29369\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__29369\,
            I => \N__29365\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__29368\,
            I => \N__29362\
        );

    \I__5174\ : Span4Mux_v
    port map (
            O => \N__29365\,
            I => \N__29359\
        );

    \I__5173\ : InMux
    port map (
            O => \N__29362\,
            I => \N__29356\
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__29359\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__29356\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__5170\ : InMux
    port map (
            O => \N__29351\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__5169\ : CascadeMux
    port map (
            O => \N__29348\,
            I => \N__29345\
        );

    \I__5168\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29342\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__29342\,
            I => \N__29339\
        );

    \I__5166\ : Span4Mux_v
    port map (
            O => \N__29339\,
            I => \N__29335\
        );

    \I__5165\ : InMux
    port map (
            O => \N__29338\,
            I => \N__29332\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__29335\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__29332\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29327\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__5161\ : InMux
    port map (
            O => \N__29324\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29321\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__5159\ : InMux
    port map (
            O => \N__29318\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__5158\ : InMux
    port map (
            O => \N__29315\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__5157\ : InMux
    port map (
            O => \N__29312\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__5156\ : InMux
    port map (
            O => \N__29309\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__5155\ : InMux
    port map (
            O => \N__29306\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__5154\ : InMux
    port map (
            O => \N__29303\,
            I => \bfn_11_17_0_\
        );

    \I__5153\ : InMux
    port map (
            O => \N__29300\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__5152\ : InMux
    port map (
            O => \N__29297\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29294\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29291\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__5149\ : InMux
    port map (
            O => \N__29288\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__5148\ : InMux
    port map (
            O => \N__29285\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__5147\ : InMux
    port map (
            O => \N__29282\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29279\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__5145\ : InMux
    port map (
            O => \N__29276\,
            I => \bfn_11_16_0_\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29268\
        );

    \I__5143\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29265\
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__29271\,
            I => \N__29260\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29268\,
            I => \N__29257\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__29265\,
            I => \N__29254\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29264\,
            I => \N__29247\
        );

    \I__5138\ : InMux
    port map (
            O => \N__29263\,
            I => \N__29247\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29260\,
            I => \N__29247\
        );

    \I__5136\ : Span4Mux_h
    port map (
            O => \N__29257\,
            I => \N__29244\
        );

    \I__5135\ : Span4Mux_h
    port map (
            O => \N__29254\,
            I => \N__29239\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__29247\,
            I => \N__29239\
        );

    \I__5133\ : Odrv4
    port map (
            O => \N__29244\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__29239\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__5131\ : InMux
    port map (
            O => \N__29234\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_31\
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__29231\,
            I => \N__29228\
        );

    \I__5129\ : InMux
    port map (
            O => \N__29228\,
            I => \N__29225\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__29225\,
            I => \N__29222\
        );

    \I__5127\ : Span4Mux_h
    port map (
            O => \N__29222\,
            I => \N__29219\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__29219\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\
        );

    \I__5125\ : CascadeMux
    port map (
            O => \N__29216\,
            I => \delay_measurement_inst.delay_hc_timer.N_382_i_cascade_\
        );

    \I__5124\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29209\
        );

    \I__5123\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29206\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__29209\,
            I => \elapsed_time_ns_1_RNIP3OD11_0_30\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__29206\,
            I => \elapsed_time_ns_1_RNIP3OD11_0_30\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__29201\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_\
        );

    \I__5119\ : CascadeMux
    port map (
            O => \N__29198\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15_cascade_\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29192\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__29192\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21\
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__29189\,
            I => \N__29185\
        );

    \I__5115\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29177\
        );

    \I__5114\ : InMux
    port map (
            O => \N__29185\,
            I => \N__29177\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29184\,
            I => \N__29177\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__29177\,
            I => \N__29174\
        );

    \I__5111\ : Odrv4
    port map (
            O => \N__29174\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\
        );

    \I__5110\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29168\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__29168\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29165\,
            I => \N__29161\
        );

    \I__5107\ : InMux
    port map (
            O => \N__29164\,
            I => \N__29158\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__29161\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__29158\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29150\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__29150\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29147\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\
        );

    \I__5101\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29141\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29138\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__29138\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\
        );

    \I__5098\ : InMux
    port map (
            O => \N__29135\,
            I => \bfn_11_13_0_\
        );

    \I__5097\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29129\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__29129\,
            I => \N__29126\
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__29126\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\
        );

    \I__5094\ : InMux
    port map (
            O => \N__29123\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__29120\,
            I => \N__29117\
        );

    \I__5092\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29114\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__29114\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\
        );

    \I__5090\ : InMux
    port map (
            O => \N__29111\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29103\
        );

    \I__5088\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29100\
        );

    \I__5087\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29097\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__29103\,
            I => \N__29092\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__29100\,
            I => \N__29092\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__29097\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__5083\ : Odrv4
    port map (
            O => \N__29092\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__5082\ : CascadeMux
    port map (
            O => \N__29087\,
            I => \N__29084\
        );

    \I__5081\ : InMux
    port map (
            O => \N__29084\,
            I => \N__29081\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__29081\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\
        );

    \I__5079\ : InMux
    port map (
            O => \N__29078\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\
        );

    \I__5078\ : InMux
    port map (
            O => \N__29075\,
            I => \N__29072\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__29072\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\
        );

    \I__5076\ : InMux
    port map (
            O => \N__29069\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\
        );

    \I__5075\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29063\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__29063\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\
        );

    \I__5073\ : InMux
    port map (
            O => \N__29060\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\
        );

    \I__5072\ : InMux
    port map (
            O => \N__29057\,
            I => \N__29053\
        );

    \I__5071\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29050\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__29053\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__29050\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__5068\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29042\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__29042\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\
        );

    \I__5066\ : InMux
    port map (
            O => \N__29039\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\
        );

    \I__5065\ : InMux
    port map (
            O => \N__29036\,
            I => \N__29032\
        );

    \I__5064\ : InMux
    port map (
            O => \N__29035\,
            I => \N__29029\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__29032\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__29029\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__5061\ : InMux
    port map (
            O => \N__29024\,
            I => \N__29021\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__29021\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\
        );

    \I__5059\ : InMux
    port map (
            O => \N__29018\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\
        );

    \I__5058\ : InMux
    port map (
            O => \N__29015\,
            I => \N__29010\
        );

    \I__5057\ : InMux
    port map (
            O => \N__29014\,
            I => \N__29007\
        );

    \I__5056\ : InMux
    port map (
            O => \N__29013\,
            I => \N__29004\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__29010\,
            I => \N__29001\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__29007\,
            I => \N__28998\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__29004\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__29001\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5051\ : Odrv12
    port map (
            O => \N__28998\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5050\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28988\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28985\
        );

    \I__5048\ : Odrv4
    port map (
            O => \N__28985\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\
        );

    \I__5047\ : InMux
    port map (
            O => \N__28982\,
            I => \bfn_11_12_0_\
        );

    \I__5046\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28976\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__28976\,
            I => \N__28971\
        );

    \I__5044\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28968\
        );

    \I__5043\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28965\
        );

    \I__5042\ : Span4Mux_h
    port map (
            O => \N__28971\,
            I => \N__28962\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__28968\,
            I => \N__28959\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__28965\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__28962\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__5038\ : Odrv12
    port map (
            O => \N__28959\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__5037\ : CascadeMux
    port map (
            O => \N__28952\,
            I => \N__28949\
        );

    \I__5036\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28946\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__28946\,
            I => \N__28943\
        );

    \I__5034\ : Odrv4
    port map (
            O => \N__28943\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\
        );

    \I__5033\ : InMux
    port map (
            O => \N__28940\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\
        );

    \I__5032\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28934\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__28934\,
            I => \N__28930\
        );

    \I__5030\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28926\
        );

    \I__5029\ : Sp12to4
    port map (
            O => \N__28930\,
            I => \N__28923\
        );

    \I__5028\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28920\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__28926\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5026\ : Odrv12
    port map (
            O => \N__28923\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__28920\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5024\ : CascadeMux
    port map (
            O => \N__28913\,
            I => \N__28910\
        );

    \I__5023\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28907\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__28907\,
            I => \N__28904\
        );

    \I__5021\ : Odrv4
    port map (
            O => \N__28904\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\
        );

    \I__5020\ : InMux
    port map (
            O => \N__28901\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\
        );

    \I__5019\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28893\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__28897\,
            I => \N__28890\
        );

    \I__5017\ : InMux
    port map (
            O => \N__28896\,
            I => \N__28887\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__28893\,
            I => \N__28884\
        );

    \I__5015\ : InMux
    port map (
            O => \N__28890\,
            I => \N__28881\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__28887\,
            I => \N__28876\
        );

    \I__5013\ : Span4Mux_v
    port map (
            O => \N__28884\,
            I => \N__28876\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__28881\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__28876\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5010\ : InMux
    port map (
            O => \N__28871\,
            I => \N__28868\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__28868\,
            I => \N__28865\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__28865\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\
        );

    \I__5007\ : InMux
    port map (
            O => \N__28862\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\
        );

    \I__5006\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28856\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__28856\,
            I => \N__28853\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__28853\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\
        );

    \I__5003\ : InMux
    port map (
            O => \N__28850\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\
        );

    \I__5002\ : CascadeMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__5001\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28841\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__28841\,
            I => \N__28836\
        );

    \I__4999\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28833\
        );

    \I__4998\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28830\
        );

    \I__4997\ : Span4Mux_h
    port map (
            O => \N__28836\,
            I => \N__28827\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__28833\,
            I => \N__28824\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__28830\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__28827\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__4993\ : Odrv12
    port map (
            O => \N__28824\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__4992\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28814\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__28814\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\
        );

    \I__4990\ : InMux
    port map (
            O => \N__28811\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\
        );

    \I__4989\ : CascadeMux
    port map (
            O => \N__28808\,
            I => \N__28805\
        );

    \I__4988\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28802\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28797\
        );

    \I__4986\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28794\
        );

    \I__4985\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28791\
        );

    \I__4984\ : Span4Mux_v
    port map (
            O => \N__28797\,
            I => \N__28788\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__28794\,
            I => \N__28785\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__28791\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__28788\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__4980\ : Odrv12
    port map (
            O => \N__28785\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__4979\ : InMux
    port map (
            O => \N__28778\,
            I => \N__28775\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__28775\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\
        );

    \I__4977\ : InMux
    port map (
            O => \N__28772\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\
        );

    \I__4976\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28766\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__28766\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_7\
        );

    \I__4974\ : InMux
    port map (
            O => \N__28763\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\
        );

    \I__4973\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28757\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__28757\,
            I => \N__28754\
        );

    \I__4971\ : Span4Mux_v
    port map (
            O => \N__28754\,
            I => \N__28751\
        );

    \I__4970\ : Span4Mux_v
    port map (
            O => \N__28751\,
            I => \N__28748\
        );

    \I__4969\ : Odrv4
    port map (
            O => \N__28748\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_8\
        );

    \I__4968\ : InMux
    port map (
            O => \N__28745\,
            I => \bfn_11_11_0_\
        );

    \I__4967\ : InMux
    port map (
            O => \N__28742\,
            I => \N__28739\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__28739\,
            I => \N__28736\
        );

    \I__4965\ : Span4Mux_h
    port map (
            O => \N__28736\,
            I => \N__28733\
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__28733\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_9\
        );

    \I__4963\ : InMux
    port map (
            O => \N__28730\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\
        );

    \I__4962\ : CascadeMux
    port map (
            O => \N__28727\,
            I => \N__28724\
        );

    \I__4961\ : InMux
    port map (
            O => \N__28724\,
            I => \N__28721\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__28721\,
            I => \N__28718\
        );

    \I__4959\ : Odrv12
    port map (
            O => \N__28718\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_10\
        );

    \I__4958\ : InMux
    port map (
            O => \N__28715\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\
        );

    \I__4957\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28709\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__28709\,
            I => \N__28706\
        );

    \I__4955\ : Span4Mux_h
    port map (
            O => \N__28706\,
            I => \N__28703\
        );

    \I__4954\ : Odrv4
    port map (
            O => \N__28703\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_11\
        );

    \I__4953\ : InMux
    port map (
            O => \N__28700\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\
        );

    \I__4952\ : InMux
    port map (
            O => \N__28697\,
            I => \N__28692\
        );

    \I__4951\ : InMux
    port map (
            O => \N__28696\,
            I => \N__28689\
        );

    \I__4950\ : InMux
    port map (
            O => \N__28695\,
            I => \N__28686\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__28692\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__28689\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__28686\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__4946\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28676\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__28676\,
            I => \N__28673\
        );

    \I__4944\ : Odrv4
    port map (
            O => \N__28673\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\
        );

    \I__4943\ : InMux
    port map (
            O => \N__28670\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\
        );

    \I__4942\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28664\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__28664\,
            I => \N__28659\
        );

    \I__4940\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28656\
        );

    \I__4939\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28653\
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__28659\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__28656\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__28653\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__4935\ : InMux
    port map (
            O => \N__28646\,
            I => \N__28643\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__28643\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\
        );

    \I__4933\ : InMux
    port map (
            O => \N__28640\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\
        );

    \I__4932\ : InMux
    port map (
            O => \N__28637\,
            I => \N__28632\
        );

    \I__4931\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28629\
        );

    \I__4930\ : InMux
    port map (
            O => \N__28635\,
            I => \N__28626\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__28632\,
            I => \N__28623\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__28629\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__28626\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__4926\ : Odrv4
    port map (
            O => \N__28623\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__28616\,
            I => \N__28613\
        );

    \I__4924\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28610\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__28610\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\
        );

    \I__4922\ : InMux
    port map (
            O => \N__28607\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__28604\,
            I => \N__28601\
        );

    \I__4920\ : InMux
    port map (
            O => \N__28601\,
            I => \N__28598\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__28598\,
            I => \N__28595\
        );

    \I__4918\ : Span4Mux_h
    port map (
            O => \N__28595\,
            I => \N__28592\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__28592\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__4916\ : CascadeMux
    port map (
            O => \N__28589\,
            I => \N__28586\
        );

    \I__4915\ : InMux
    port map (
            O => \N__28586\,
            I => \N__28583\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__28583\,
            I => \N__28580\
        );

    \I__4913\ : Span4Mux_h
    port map (
            O => \N__28580\,
            I => \N__28577\
        );

    \I__4912\ : Odrv4
    port map (
            O => \N__28577\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__4911\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28570\
        );

    \I__4910\ : InMux
    port map (
            O => \N__28573\,
            I => \N__28567\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__28570\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__28567\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__4907\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28559\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__28559\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\
        );

    \I__4905\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28553\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__28553\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\
        );

    \I__4903\ : InMux
    port map (
            O => \N__28550\,
            I => \N__28547\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__28547\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\
        );

    \I__4901\ : InMux
    port map (
            O => \N__28544\,
            I => \N__28541\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__28541\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\
        );

    \I__4899\ : InMux
    port map (
            O => \N__28538\,
            I => \N__28535\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__28535\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_4\
        );

    \I__4897\ : InMux
    port map (
            O => \N__28532\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\
        );

    \I__4896\ : CascadeMux
    port map (
            O => \N__28529\,
            I => \N__28526\
        );

    \I__4895\ : InMux
    port map (
            O => \N__28526\,
            I => \N__28523\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__28523\,
            I => \N__28520\
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__28520\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_5\
        );

    \I__4892\ : InMux
    port map (
            O => \N__28517\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\
        );

    \I__4891\ : InMux
    port map (
            O => \N__28514\,
            I => \N__28511\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__28511\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_6\
        );

    \I__4889\ : InMux
    port map (
            O => \N__28508\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\
        );

    \I__4888\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28502\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__28502\,
            I => \N__28499\
        );

    \I__4886\ : Span4Mux_h
    port map (
            O => \N__28499\,
            I => \N__28496\
        );

    \I__4885\ : Span4Mux_h
    port map (
            O => \N__28496\,
            I => \N__28493\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__28493\,
            I => \current_shift_inst.PI_CTRL.integrator_i_19\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__28490\,
            I => \N__28487\
        );

    \I__4882\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28484\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__28484\,
            I => \N__28480\
        );

    \I__4880\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28475\
        );

    \I__4879\ : Span4Mux_v
    port map (
            O => \N__28480\,
            I => \N__28472\
        );

    \I__4878\ : CascadeMux
    port map (
            O => \N__28479\,
            I => \N__28469\
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__28478\,
            I => \N__28466\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__28475\,
            I => \N__28462\
        );

    \I__4875\ : Span4Mux_h
    port map (
            O => \N__28472\,
            I => \N__28459\
        );

    \I__4874\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28454\
        );

    \I__4873\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28454\
        );

    \I__4872\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28451\
        );

    \I__4871\ : Odrv4
    port map (
            O => \N__28462\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4870\ : Odrv4
    port map (
            O => \N__28459\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__28454\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__28451\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__28442\,
            I => \N__28439\
        );

    \I__4866\ : InMux
    port map (
            O => \N__28439\,
            I => \N__28436\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__28436\,
            I => \N__28433\
        );

    \I__4864\ : Span4Mux_v
    port map (
            O => \N__28433\,
            I => \N__28430\
        );

    \I__4863\ : Odrv4
    port map (
            O => \N__28430\,
            I => \current_shift_inst.PI_CTRL.integrator_i_12\
        );

    \I__4862\ : InMux
    port map (
            O => \N__28427\,
            I => \N__28423\
        );

    \I__4861\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28420\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__28423\,
            I => \N__28416\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__28420\,
            I => \N__28412\
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__28419\,
            I => \N__28409\
        );

    \I__4857\ : Span4Mux_v
    port map (
            O => \N__28416\,
            I => \N__28405\
        );

    \I__4856\ : InMux
    port map (
            O => \N__28415\,
            I => \N__28402\
        );

    \I__4855\ : Span4Mux_h
    port map (
            O => \N__28412\,
            I => \N__28399\
        );

    \I__4854\ : InMux
    port map (
            O => \N__28409\,
            I => \N__28396\
        );

    \I__4853\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28393\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__28405\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__28402\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__28399\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__28396\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__28393\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4847\ : CascadeMux
    port map (
            O => \N__28382\,
            I => \N__28379\
        );

    \I__4846\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28376\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__28376\,
            I => \N__28373\
        );

    \I__4844\ : Odrv4
    port map (
            O => \N__28373\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__28370\,
            I => \N__28367\
        );

    \I__4842\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28364\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__28364\,
            I => \N__28361\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__28361\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\
        );

    \I__4839\ : InMux
    port map (
            O => \N__28358\,
            I => \N__28355\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__28355\,
            I => \N__28352\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__28352\,
            I => \N__28349\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__28349\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__4835\ : InMux
    port map (
            O => \N__28346\,
            I => \N__28343\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__28343\,
            I => \N__28340\
        );

    \I__4833\ : Odrv12
    port map (
            O => \N__28340\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__4832\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28334\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__28334\,
            I => \N__28331\
        );

    \I__4830\ : Odrv12
    port map (
            O => \N__28331\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__4829\ : InMux
    port map (
            O => \N__28328\,
            I => \N__28325\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__28325\,
            I => \N__28322\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__28322\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__28319\,
            I => \N__28310\
        );

    \I__4825\ : InMux
    port map (
            O => \N__28318\,
            I => \N__28293\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28317\,
            I => \N__28290\
        );

    \I__4823\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28281\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28315\,
            I => \N__28281\
        );

    \I__4821\ : InMux
    port map (
            O => \N__28314\,
            I => \N__28281\
        );

    \I__4820\ : InMux
    port map (
            O => \N__28313\,
            I => \N__28281\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28270\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28270\
        );

    \I__4817\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28270\
        );

    \I__4816\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28270\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28270\
        );

    \I__4814\ : InMux
    port map (
            O => \N__28305\,
            I => \N__28257\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28246\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28303\,
            I => \N__28246\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28246\
        );

    \I__4810\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28246\
        );

    \I__4809\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28246\
        );

    \I__4808\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28237\
        );

    \I__4807\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28237\
        );

    \I__4806\ : InMux
    port map (
            O => \N__28297\,
            I => \N__28237\
        );

    \I__4805\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28237\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__28293\,
            I => \N__28234\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__28290\,
            I => \N__28230\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__28281\,
            I => \N__28225\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__28270\,
            I => \N__28225\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28222\
        );

    \I__4799\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28211\
        );

    \I__4798\ : InMux
    port map (
            O => \N__28267\,
            I => \N__28211\
        );

    \I__4797\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28211\
        );

    \I__4796\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28211\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28211\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28263\,
            I => \N__28202\
        );

    \I__4793\ : InMux
    port map (
            O => \N__28262\,
            I => \N__28202\
        );

    \I__4792\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28202\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28202\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__28257\,
            I => \N__28199\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__28246\,
            I => \N__28194\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__28237\,
            I => \N__28194\
        );

    \I__4787\ : Span4Mux_v
    port map (
            O => \N__28234\,
            I => \N__28191\
        );

    \I__4786\ : InMux
    port map (
            O => \N__28233\,
            I => \N__28188\
        );

    \I__4785\ : Span4Mux_h
    port map (
            O => \N__28230\,
            I => \N__28183\
        );

    \I__4784\ : Span4Mux_h
    port map (
            O => \N__28225\,
            I => \N__28183\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__28222\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__28211\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__28202\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__28199\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4779\ : Odrv4
    port map (
            O => \N__28194\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__28191\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__28188\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__28183\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4775\ : CascadeMux
    port map (
            O => \N__28166\,
            I => \N__28153\
        );

    \I__4774\ : CascadeMux
    port map (
            O => \N__28165\,
            I => \N__28140\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__28164\,
            I => \N__28136\
        );

    \I__4772\ : CascadeMux
    port map (
            O => \N__28163\,
            I => \N__28133\
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__28162\,
            I => \N__28130\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__28161\,
            I => \N__28126\
        );

    \I__4769\ : CascadeMux
    port map (
            O => \N__28160\,
            I => \N__28123\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28114\
        );

    \I__4767\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28114\
        );

    \I__4766\ : InMux
    port map (
            O => \N__28157\,
            I => \N__28114\
        );

    \I__4765\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28114\
        );

    \I__4764\ : InMux
    port map (
            O => \N__28153\,
            I => \N__28111\
        );

    \I__4763\ : CascadeMux
    port map (
            O => \N__28152\,
            I => \N__28108\
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__28151\,
            I => \N__28105\
        );

    \I__4761\ : CascadeMux
    port map (
            O => \N__28150\,
            I => \N__28102\
        );

    \I__4760\ : CascadeMux
    port map (
            O => \N__28149\,
            I => \N__28095\
        );

    \I__4759\ : CascadeMux
    port map (
            O => \N__28148\,
            I => \N__28092\
        );

    \I__4758\ : CascadeMux
    port map (
            O => \N__28147\,
            I => \N__28089\
        );

    \I__4757\ : CascadeMux
    port map (
            O => \N__28146\,
            I => \N__28086\
        );

    \I__4756\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28077\
        );

    \I__4755\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28077\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28077\
        );

    \I__4753\ : InMux
    port map (
            O => \N__28140\,
            I => \N__28077\
        );

    \I__4752\ : InMux
    port map (
            O => \N__28139\,
            I => \N__28068\
        );

    \I__4751\ : InMux
    port map (
            O => \N__28136\,
            I => \N__28068\
        );

    \I__4750\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28068\
        );

    \I__4749\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28068\
        );

    \I__4748\ : InMux
    port map (
            O => \N__28129\,
            I => \N__28061\
        );

    \I__4747\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28061\
        );

    \I__4746\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28061\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28114\,
            I => \N__28056\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__28111\,
            I => \N__28056\
        );

    \I__4743\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28053\
        );

    \I__4742\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28046\
        );

    \I__4741\ : InMux
    port map (
            O => \N__28102\,
            I => \N__28046\
        );

    \I__4740\ : InMux
    port map (
            O => \N__28101\,
            I => \N__28046\
        );

    \I__4739\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28035\
        );

    \I__4738\ : InMux
    port map (
            O => \N__28099\,
            I => \N__28035\
        );

    \I__4737\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28035\
        );

    \I__4736\ : InMux
    port map (
            O => \N__28095\,
            I => \N__28035\
        );

    \I__4735\ : InMux
    port map (
            O => \N__28092\,
            I => \N__28035\
        );

    \I__4734\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28030\
        );

    \I__4733\ : InMux
    port map (
            O => \N__28086\,
            I => \N__28030\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__28077\,
            I => \N__28027\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__28068\,
            I => \N__28024\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__28061\,
            I => \N__28019\
        );

    \I__4729\ : Span4Mux_v
    port map (
            O => \N__28056\,
            I => \N__28019\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__28053\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__28046\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__28035\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__28030\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4724\ : Odrv4
    port map (
            O => \N__28027\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4723\ : Odrv4
    port map (
            O => \N__28024\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__28019\,
            I => \current_shift_inst.PI_CTRL.N_103\
        );

    \I__4721\ : InMux
    port map (
            O => \N__28004\,
            I => \N__27985\
        );

    \I__4720\ : InMux
    port map (
            O => \N__28003\,
            I => \N__27985\
        );

    \I__4719\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27985\
        );

    \I__4718\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27985\
        );

    \I__4717\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27985\
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__27999\,
            I => \N__27971\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__27998\,
            I => \N__27968\
        );

    \I__4714\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27962\
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__27996\,
            I => \N__27957\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__27985\,
            I => \N__27948\
        );

    \I__4711\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27939\
        );

    \I__4710\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27939\
        );

    \I__4709\ : InMux
    port map (
            O => \N__27982\,
            I => \N__27939\
        );

    \I__4708\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27939\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__27980\,
            I => \N__27936\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__27979\,
            I => \N__27932\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__27978\,
            I => \N__27929\
        );

    \I__4704\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27926\
        );

    \I__4703\ : InMux
    port map (
            O => \N__27976\,
            I => \N__27921\
        );

    \I__4702\ : InMux
    port map (
            O => \N__27975\,
            I => \N__27921\
        );

    \I__4701\ : InMux
    port map (
            O => \N__27974\,
            I => \N__27912\
        );

    \I__4700\ : InMux
    port map (
            O => \N__27971\,
            I => \N__27912\
        );

    \I__4699\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27912\
        );

    \I__4698\ : InMux
    port map (
            O => \N__27967\,
            I => \N__27912\
        );

    \I__4697\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27907\
        );

    \I__4696\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27907\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__27962\,
            I => \N__27904\
        );

    \I__4694\ : InMux
    port map (
            O => \N__27961\,
            I => \N__27901\
        );

    \I__4693\ : InMux
    port map (
            O => \N__27960\,
            I => \N__27892\
        );

    \I__4692\ : InMux
    port map (
            O => \N__27957\,
            I => \N__27892\
        );

    \I__4691\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27892\
        );

    \I__4690\ : InMux
    port map (
            O => \N__27955\,
            I => \N__27892\
        );

    \I__4689\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27883\
        );

    \I__4688\ : InMux
    port map (
            O => \N__27953\,
            I => \N__27883\
        );

    \I__4687\ : InMux
    port map (
            O => \N__27952\,
            I => \N__27883\
        );

    \I__4686\ : InMux
    port map (
            O => \N__27951\,
            I => \N__27883\
        );

    \I__4685\ : Span4Mux_v
    port map (
            O => \N__27948\,
            I => \N__27878\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__27939\,
            I => \N__27878\
        );

    \I__4683\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27875\
        );

    \I__4682\ : InMux
    port map (
            O => \N__27935\,
            I => \N__27868\
        );

    \I__4681\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27868\
        );

    \I__4680\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27868\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27865\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__27921\,
            I => \N__27856\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__27912\,
            I => \N__27856\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__27907\,
            I => \N__27856\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__27904\,
            I => \N__27856\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__27901\,
            I => \N__27847\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__27892\,
            I => \N__27847\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__27883\,
            I => \N__27847\
        );

    \I__4671\ : Span4Mux_v
    port map (
            O => \N__27878\,
            I => \N__27847\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__27875\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__27868\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4668\ : Odrv4
    port map (
            O => \N__27865\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4667\ : Odrv4
    port map (
            O => \N__27856\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4666\ : Odrv4
    port map (
            O => \N__27847\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__27836\,
            I => \N__27833\
        );

    \I__4664\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27828\
        );

    \I__4663\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27825\
        );

    \I__4662\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27822\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__27828\,
            I => \N__27810\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__27825\,
            I => \N__27810\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__27822\,
            I => \N__27810\
        );

    \I__4658\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27805\
        );

    \I__4657\ : InMux
    port map (
            O => \N__27820\,
            I => \N__27805\
        );

    \I__4656\ : InMux
    port map (
            O => \N__27819\,
            I => \N__27802\
        );

    \I__4655\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27799\
        );

    \I__4654\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27796\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__27810\,
            I => \N__27793\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__27805\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__27802\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__27799\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__27796\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__27793\,
            I => \elapsed_time_ns_1_RNIS4MD11_0_15\
        );

    \I__4647\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27778\
        );

    \I__4646\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27775\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__27778\,
            I => \N__27772\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__27775\,
            I => \N__27769\
        );

    \I__4643\ : Span4Mux_v
    port map (
            O => \N__27772\,
            I => \N__27766\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__27769\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__27766\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO\
        );

    \I__4640\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27758\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__27758\,
            I => \N__27755\
        );

    \I__4638\ : Odrv12
    port map (
            O => \N__27755\,
            I => \phase_controller_inst2.stoper_hc.running_1_sqmuxa\
        );

    \I__4637\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27744\
        );

    \I__4636\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27744\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__27750\,
            I => \N__27740\
        );

    \I__4634\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27735\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__27744\,
            I => \N__27732\
        );

    \I__4632\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27725\
        );

    \I__4631\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27725\
        );

    \I__4630\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27725\
        );

    \I__4629\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27722\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27719\
        );

    \I__4627\ : Span4Mux_h
    port map (
            O => \N__27732\,
            I => \N__27714\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__27725\,
            I => \N__27714\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__27722\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__4624\ : Odrv12
    port map (
            O => \N__27719\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__27714\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__4622\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27700\
        );

    \I__4621\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27700\
        );

    \I__4620\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27693\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__27700\,
            I => \N__27690\
        );

    \I__4618\ : InMux
    port map (
            O => \N__27699\,
            I => \N__27681\
        );

    \I__4617\ : InMux
    port map (
            O => \N__27698\,
            I => \N__27681\
        );

    \I__4616\ : InMux
    port map (
            O => \N__27697\,
            I => \N__27681\
        );

    \I__4615\ : InMux
    port map (
            O => \N__27696\,
            I => \N__27681\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__27693\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__27690\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__27681\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4611\ : CascadeMux
    port map (
            O => \N__27674\,
            I => \phase_controller_inst2.stoper_hc.running_1_sqmuxa_cascade_\
        );

    \I__4610\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27668\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__27668\,
            I => \N__27663\
        );

    \I__4608\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27658\
        );

    \I__4607\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27658\
        );

    \I__4606\ : Odrv4
    port map (
            O => \N__27663\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__27658\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__4604\ : InMux
    port map (
            O => \N__27653\,
            I => \N__27650\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__27650\,
            I => \N__27647\
        );

    \I__4602\ : Odrv12
    port map (
            O => \N__27647\,
            I => \phase_controller_inst2.stoper_hc.un1_start_latched2_0\
        );

    \I__4601\ : IoInMux
    port map (
            O => \N__27644\,
            I => \N__27641\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__27641\,
            I => \N__27638\
        );

    \I__4599\ : Span4Mux_s2_v
    port map (
            O => \N__27638\,
            I => \N__27635\
        );

    \I__4598\ : Span4Mux_v
    port map (
            O => \N__27635\,
            I => \N__27632\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__27632\,
            I => s4_phy_c
        );

    \I__4596\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27626\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__27626\,
            I => \N__27623\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__27623\,
            I => \il_max_comp1_D1\
        );

    \I__4593\ : InMux
    port map (
            O => \N__27620\,
            I => \N__27617\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__27617\,
            I => \N__27614\
        );

    \I__4591\ : Span4Mux_v
    port map (
            O => \N__27614\,
            I => \N__27611\
        );

    \I__4590\ : Span4Mux_h
    port map (
            O => \N__27611\,
            I => \N__27608\
        );

    \I__4589\ : Odrv4
    port map (
            O => \N__27608\,
            I => il_min_comp2_c
        );

    \I__4588\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27602\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__27602\,
            I => \il_min_comp2_D1\
        );

    \I__4586\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27592\
        );

    \I__4585\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27589\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__27597\,
            I => \N__27586\
        );

    \I__4583\ : CascadeMux
    port map (
            O => \N__27596\,
            I => \N__27583\
        );

    \I__4582\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27580\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__27592\,
            I => \N__27577\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__27589\,
            I => \N__27574\
        );

    \I__4579\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27571\
        );

    \I__4578\ : InMux
    port map (
            O => \N__27583\,
            I => \N__27568\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__27580\,
            I => \N__27565\
        );

    \I__4576\ : Span4Mux_v
    port map (
            O => \N__27577\,
            I => \N__27562\
        );

    \I__4575\ : Span4Mux_v
    port map (
            O => \N__27574\,
            I => \N__27555\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__27571\,
            I => \N__27555\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__27568\,
            I => \N__27555\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__27565\,
            I => \N__27552\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__27562\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__27555\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__4569\ : Odrv4
    port map (
            O => \N__27552\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__4568\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__27542\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5\
        );

    \I__4566\ : CascadeMux
    port map (
            O => \N__27539\,
            I => \N__27536\
        );

    \I__4565\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27533\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__27533\,
            I => \N__27530\
        );

    \I__4563\ : Span4Mux_h
    port map (
            O => \N__27530\,
            I => \N__27526\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27522\
        );

    \I__4561\ : Span4Mux_h
    port map (
            O => \N__27526\,
            I => \N__27519\
        );

    \I__4560\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27516\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__27522\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__27519\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__27516\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10\
        );

    \I__4556\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27506\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__27506\,
            I => \N__27500\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__27505\,
            I => \N__27497\
        );

    \I__4553\ : InMux
    port map (
            O => \N__27504\,
            I => \N__27494\
        );

    \I__4552\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27491\
        );

    \I__4551\ : Span4Mux_h
    port map (
            O => \N__27500\,
            I => \N__27488\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27485\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__27494\,
            I => \N__27482\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__27491\,
            I => \elapsed_time_ns_1_RNIQ2MD11_0_13\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__27488\,
            I => \elapsed_time_ns_1_RNIQ2MD11_0_13\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__27485\,
            I => \elapsed_time_ns_1_RNIQ2MD11_0_13\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__27482\,
            I => \elapsed_time_ns_1_RNIQ2MD11_0_13\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__27473\,
            I => \elapsed_time_ns_1_RNINVLD11_0_10_cascade_\
        );

    \I__4543\ : CascadeMux
    port map (
            O => \N__27470\,
            I => \N__27466\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__27469\,
            I => \N__27463\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27460\
        );

    \I__4540\ : InMux
    port map (
            O => \N__27463\,
            I => \N__27457\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__27460\,
            I => \N__27454\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__27457\,
            I => \N__27449\
        );

    \I__4537\ : Span4Mux_h
    port map (
            O => \N__27454\,
            I => \N__27449\
        );

    \I__4536\ : Span4Mux_h
    port map (
            O => \N__27449\,
            I => \N__27444\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27439\
        );

    \I__4534\ : InMux
    port map (
            O => \N__27447\,
            I => \N__27439\
        );

    \I__4533\ : Odrv4
    port map (
            O => \N__27444\,
            I => \elapsed_time_ns_1_RNIP1MD11_0_12\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__27439\,
            I => \elapsed_time_ns_1_RNIP1MD11_0_12\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__27434\,
            I => \phase_controller_inst1.stoper_hc.N_319_cascade_\
        );

    \I__4530\ : CascadeMux
    port map (
            O => \N__27431\,
            I => \N__27428\
        );

    \I__4529\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27423\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27420\
        );

    \I__4527\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27417\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__27423\,
            I => \N__27413\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__27420\,
            I => \N__27408\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__27417\,
            I => \N__27408\
        );

    \I__4523\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27405\
        );

    \I__4522\ : Span12Mux_s10_h
    port map (
            O => \N__27413\,
            I => \N__27400\
        );

    \I__4521\ : Sp12to4
    port map (
            O => \N__27408\,
            I => \N__27395\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__27405\,
            I => \N__27395\
        );

    \I__4519\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27390\
        );

    \I__4518\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27390\
        );

    \I__4517\ : Odrv12
    port map (
            O => \N__27400\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__4516\ : Odrv12
    port map (
            O => \N__27395\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__27390\,
            I => \elapsed_time_ns_1_RNI1TBED1_0_14\
        );

    \I__4514\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27380\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__27380\,
            I => \phase_controller_inst1.stoper_hc.N_275\
        );

    \I__4512\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27373\
        );

    \I__4511\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27370\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__27373\,
            I => \phase_controller_inst1.stoper_hc.N_319\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__27370\,
            I => \phase_controller_inst1.stoper_hc.N_319\
        );

    \I__4508\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27362\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__27362\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0Z0Z_9\
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__27359\,
            I => \N__27351\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27358\,
            I => \N__27333\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27326\
        );

    \I__4503\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27326\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27326\
        );

    \I__4501\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27315\
        );

    \I__4500\ : InMux
    port map (
            O => \N__27351\,
            I => \N__27315\
        );

    \I__4499\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27315\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27315\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27315\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27306\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27306\
        );

    \I__4494\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27306\
        );

    \I__4493\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27306\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__27343\,
            I => \N__27301\
        );

    \I__4491\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27277\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27277\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27277\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27277\
        );

    \I__4487\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27277\
        );

    \I__4486\ : InMux
    port map (
            O => \N__27337\,
            I => \N__27277\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27277\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27333\,
            I => \N__27270\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__27326\,
            I => \N__27270\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__27315\,
            I => \N__27270\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__27306\,
            I => \N__27267\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27263\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27256\
        );

    \I__4478\ : InMux
    port map (
            O => \N__27301\,
            I => \N__27256\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27300\,
            I => \N__27256\
        );

    \I__4476\ : CascadeMux
    port map (
            O => \N__27299\,
            I => \N__27252\
        );

    \I__4475\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27248\
        );

    \I__4474\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27235\
        );

    \I__4473\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27235\
        );

    \I__4472\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27235\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27235\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27235\
        );

    \I__4469\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27235\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__27277\,
            I => \N__27232\
        );

    \I__4467\ : Sp12to4
    port map (
            O => \N__27270\,
            I => \N__27227\
        );

    \I__4466\ : Span12Mux_s9_h
    port map (
            O => \N__27267\,
            I => \N__27227\
        );

    \I__4465\ : InMux
    port map (
            O => \N__27266\,
            I => \N__27224\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__27263\,
            I => \N__27219\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__27256\,
            I => \N__27219\
        );

    \I__4462\ : InMux
    port map (
            O => \N__27255\,
            I => \N__27212\
        );

    \I__4461\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27212\
        );

    \I__4460\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27212\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__27248\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__27235\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__27232\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4456\ : Odrv12
    port map (
            O => \N__27227\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__27224\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__27219\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__27212\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__27197\,
            I => \N__27193\
        );

    \I__4451\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27189\
        );

    \I__4450\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27185\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27192\,
            I => \N__27182\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__27189\,
            I => \N__27179\
        );

    \I__4447\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27176\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__27185\,
            I => \N__27171\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__27182\,
            I => \N__27171\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__27179\,
            I => \phase_controller_inst1.stoper_hc.N_278\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__27176\,
            I => \phase_controller_inst1.stoper_hc.N_278\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__27171\,
            I => \phase_controller_inst1.stoper_hc.N_278\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27164\,
            I => \N__27151\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27151\
        );

    \I__4439\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27151\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27151\
        );

    \I__4437\ : CascadeMux
    port map (
            O => \N__27160\,
            I => \N__27143\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__27151\,
            I => \N__27139\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27150\,
            I => \N__27136\
        );

    \I__4434\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27133\
        );

    \I__4433\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27126\
        );

    \I__4432\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27126\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27126\
        );

    \I__4430\ : InMux
    port map (
            O => \N__27143\,
            I => \N__27123\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27142\,
            I => \N__27107\
        );

    \I__4428\ : Span4Mux_h
    port map (
            O => \N__27139\,
            I => \N__27102\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__27136\,
            I => \N__27093\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__27133\,
            I => \N__27093\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__27126\,
            I => \N__27093\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__27123\,
            I => \N__27093\
        );

    \I__4423\ : InMux
    port map (
            O => \N__27122\,
            I => \N__27090\
        );

    \I__4422\ : InMux
    port map (
            O => \N__27121\,
            I => \N__27085\
        );

    \I__4421\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27085\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27076\
        );

    \I__4419\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27076\
        );

    \I__4418\ : InMux
    port map (
            O => \N__27117\,
            I => \N__27076\
        );

    \I__4417\ : InMux
    port map (
            O => \N__27116\,
            I => \N__27076\
        );

    \I__4416\ : InMux
    port map (
            O => \N__27115\,
            I => \N__27063\
        );

    \I__4415\ : InMux
    port map (
            O => \N__27114\,
            I => \N__27063\
        );

    \I__4414\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27063\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27063\
        );

    \I__4412\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27063\
        );

    \I__4411\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27063\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27060\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27106\,
            I => \N__27055\
        );

    \I__4408\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27055\
        );

    \I__4407\ : Span4Mux_h
    port map (
            O => \N__27102\,
            I => \N__27050\
        );

    \I__4406\ : Span4Mux_v
    port map (
            O => \N__27093\,
            I => \N__27050\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__27090\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__27085\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__27076\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__27063\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4401\ : Odrv12
    port map (
            O => \N__27060\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__27055\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__27050\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__27035\,
            I => \N__27032\
        );

    \I__4397\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__27029\,
            I => \N__27026\
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__27026\,
            I => \phase_controller_inst2.stoper_hc.un6_running_15\
        );

    \I__4394\ : CEMux
    port map (
            O => \N__27023\,
            I => \N__27017\
        );

    \I__4393\ : CEMux
    port map (
            O => \N__27022\,
            I => \N__27010\
        );

    \I__4392\ : CEMux
    port map (
            O => \N__27021\,
            I => \N__27003\
        );

    \I__4391\ : CEMux
    port map (
            O => \N__27020\,
            I => \N__27000\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__27017\,
            I => \N__26997\
        );

    \I__4389\ : CEMux
    port map (
            O => \N__27016\,
            I => \N__26994\
        );

    \I__4388\ : InMux
    port map (
            O => \N__27015\,
            I => \N__26991\
        );

    \I__4387\ : CEMux
    port map (
            O => \N__27014\,
            I => \N__26988\
        );

    \I__4386\ : CEMux
    port map (
            O => \N__27013\,
            I => \N__26985\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__27010\,
            I => \N__26982\
        );

    \I__4384\ : InMux
    port map (
            O => \N__27009\,
            I => \N__26973\
        );

    \I__4383\ : InMux
    port map (
            O => \N__27008\,
            I => \N__26973\
        );

    \I__4382\ : InMux
    port map (
            O => \N__27007\,
            I => \N__26973\
        );

    \I__4381\ : InMux
    port map (
            O => \N__27006\,
            I => \N__26973\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__27003\,
            I => \N__26970\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__27000\,
            I => \N__26967\
        );

    \I__4378\ : Span4Mux_h
    port map (
            O => \N__26997\,
            I => \N__26950\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__26994\,
            I => \N__26947\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__26991\,
            I => \N__26942\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__26988\,
            I => \N__26942\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__26985\,
            I => \N__26939\
        );

    \I__4373\ : Span4Mux_h
    port map (
            O => \N__26982\,
            I => \N__26936\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__26973\,
            I => \N__26929\
        );

    \I__4371\ : Span4Mux_v
    port map (
            O => \N__26970\,
            I => \N__26929\
        );

    \I__4370\ : Span4Mux_v
    port map (
            O => \N__26967\,
            I => \N__26929\
        );

    \I__4369\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26922\
        );

    \I__4368\ : InMux
    port map (
            O => \N__26965\,
            I => \N__26922\
        );

    \I__4367\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26922\
        );

    \I__4366\ : InMux
    port map (
            O => \N__26963\,
            I => \N__26913\
        );

    \I__4365\ : InMux
    port map (
            O => \N__26962\,
            I => \N__26913\
        );

    \I__4364\ : InMux
    port map (
            O => \N__26961\,
            I => \N__26913\
        );

    \I__4363\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26913\
        );

    \I__4362\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26910\
        );

    \I__4361\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26905\
        );

    \I__4360\ : InMux
    port map (
            O => \N__26957\,
            I => \N__26905\
        );

    \I__4359\ : InMux
    port map (
            O => \N__26956\,
            I => \N__26896\
        );

    \I__4358\ : InMux
    port map (
            O => \N__26955\,
            I => \N__26896\
        );

    \I__4357\ : InMux
    port map (
            O => \N__26954\,
            I => \N__26896\
        );

    \I__4356\ : InMux
    port map (
            O => \N__26953\,
            I => \N__26896\
        );

    \I__4355\ : Span4Mux_v
    port map (
            O => \N__26950\,
            I => \N__26893\
        );

    \I__4354\ : Span4Mux_h
    port map (
            O => \N__26947\,
            I => \N__26888\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__26942\,
            I => \N__26888\
        );

    \I__4352\ : Span12Mux_v
    port map (
            O => \N__26939\,
            I => \N__26885\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__26936\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4350\ : Odrv4
    port map (
            O => \N__26929\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__26922\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__26913\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__26910\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__26905\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__26896\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__26893\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__26888\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4342\ : Odrv12
    port map (
            O => \N__26885\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4341\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26861\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__26861\,
            I => \N__26857\
        );

    \I__4339\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26854\
        );

    \I__4338\ : Span4Mux_h
    port map (
            O => \N__26857\,
            I => \N__26848\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__26854\,
            I => \N__26848\
        );

    \I__4336\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26844\
        );

    \I__4335\ : Span4Mux_v
    port map (
            O => \N__26848\,
            I => \N__26841\
        );

    \I__4334\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26838\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__26844\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__26841\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__26838\,
            I => \elapsed_time_ns_1_RNID6DJ11_0_7\
        );

    \I__4330\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26828\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__26828\,
            I => \N__26823\
        );

    \I__4328\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26820\
        );

    \I__4327\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26816\
        );

    \I__4326\ : Span4Mux_h
    port map (
            O => \N__26823\,
            I => \N__26813\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26810\
        );

    \I__4324\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26807\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__26816\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__26813\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__26810\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__26807\,
            I => \elapsed_time_ns_1_RNIE7DJ11_0_8\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__26798\,
            I => \N__26794\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__26797\,
            I => \N__26791\
        );

    \I__4317\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26788\
        );

    \I__4316\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26783\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__26788\,
            I => \N__26780\
        );

    \I__4314\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26777\
        );

    \I__4313\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26774\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__26783\,
            I => \N__26771\
        );

    \I__4311\ : Span4Mux_h
    port map (
            O => \N__26780\,
            I => \N__26768\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__26777\,
            I => \N__26765\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__26774\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__26771\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__26768\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__26765\,
            I => \elapsed_time_ns_1_RNIB4DJ11_0_5\
        );

    \I__4305\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26753\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__26753\,
            I => \N__26745\
        );

    \I__4303\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26742\
        );

    \I__4302\ : InMux
    port map (
            O => \N__26751\,
            I => \N__26739\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26736\
        );

    \I__4300\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26731\
        );

    \I__4299\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26728\
        );

    \I__4298\ : Span4Mux_v
    port map (
            O => \N__26745\,
            I => \N__26719\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__26742\,
            I => \N__26719\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__26739\,
            I => \N__26719\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__26736\,
            I => \N__26719\
        );

    \I__4294\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26714\
        );

    \I__4293\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26714\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__26731\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__26728\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__4290\ : Odrv4
    port map (
            O => \N__26719\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__26714\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__26705\,
            I => \elapsed_time_ns_1_RNI3VBED1_0_16_cascade_\
        );

    \I__4287\ : InMux
    port map (
            O => \N__26702\,
            I => \N__26699\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26695\
        );

    \I__4285\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26692\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__26695\,
            I => \N__26688\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__26692\,
            I => \N__26685\
        );

    \I__4282\ : InMux
    port map (
            O => \N__26691\,
            I => \N__26682\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__26688\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4280\ : Odrv4
    port map (
            O => \N__26685\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__26682\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4\
        );

    \I__4278\ : InMux
    port map (
            O => \N__26675\,
            I => \N__26668\
        );

    \I__4277\ : InMux
    port map (
            O => \N__26674\,
            I => \N__26663\
        );

    \I__4276\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26663\
        );

    \I__4275\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26658\
        );

    \I__4274\ : InMux
    port map (
            O => \N__26671\,
            I => \N__26658\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__26668\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__26663\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__26658\,
            I => \elapsed_time_ns_1_RNI40CED1_0_17\
        );

    \I__4270\ : CascadeMux
    port map (
            O => \N__26651\,
            I => \elapsed_time_ns_1_RNIA3DJ11_0_4_cascade_\
        );

    \I__4269\ : InMux
    port map (
            O => \N__26648\,
            I => \N__26643\
        );

    \I__4268\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26640\
        );

    \I__4267\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26635\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__26643\,
            I => \N__26630\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__26640\,
            I => \N__26630\
        );

    \I__4264\ : InMux
    port map (
            O => \N__26639\,
            I => \N__26625\
        );

    \I__4263\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26625\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__26635\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__4261\ : Odrv12
    port map (
            O => \N__26630\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__26625\,
            I => \elapsed_time_ns_1_RNI51CED1_0_18\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__26618\,
            I => \N__26614\
        );

    \I__4258\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26609\
        );

    \I__4257\ : InMux
    port map (
            O => \N__26614\,
            I => \N__26604\
        );

    \I__4256\ : InMux
    port map (
            O => \N__26613\,
            I => \N__26604\
        );

    \I__4255\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26601\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__26609\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__26604\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__26601\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__26594\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_\
        );

    \I__4250\ : InMux
    port map (
            O => \N__26591\,
            I => \N__26587\
        );

    \I__4249\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26584\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__26587\,
            I => \N__26579\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__26584\,
            I => \N__26579\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__26579\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__4245\ : CascadeMux
    port map (
            O => \N__26576\,
            I => \N__26571\
        );

    \I__4244\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26564\
        );

    \I__4243\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26564\
        );

    \I__4242\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26564\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__26564\,
            I => \phase_controller_inst1.stoper_hc.N_337\
        );

    \I__4240\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26558\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__26558\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4\
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__26555\,
            I => \N__26551\
        );

    \I__4237\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26547\
        );

    \I__4236\ : InMux
    port map (
            O => \N__26551\,
            I => \N__26544\
        );

    \I__4235\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26541\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__26547\,
            I => \N__26538\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__26544\,
            I => \N__26533\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__26541\,
            I => \N__26528\
        );

    \I__4231\ : Span4Mux_v
    port map (
            O => \N__26538\,
            I => \N__26528\
        );

    \I__4230\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26523\
        );

    \I__4229\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26523\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__26533\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__26528\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__26523\,
            I => \elapsed_time_ns_1_RNIQURR91_0_3\
        );

    \I__4225\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26513\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__26513\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__26510\,
            I => \N__26507\
        );

    \I__4222\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26503\
        );

    \I__4221\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26500\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26497\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__26500\,
            I => \elapsed_time_ns_1_RNIP2ND11_0_21\
        );

    \I__4218\ : Odrv12
    port map (
            O => \N__26497\,
            I => \elapsed_time_ns_1_RNIP2ND11_0_21\
        );

    \I__4217\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26488\
        );

    \I__4216\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26485\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__26488\,
            I => \elapsed_time_ns_1_RNIS5ND11_0_24\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__26485\,
            I => \elapsed_time_ns_1_RNIS5ND11_0_24\
        );

    \I__4213\ : InMux
    port map (
            O => \N__26480\,
            I => \N__26477\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__26477\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__26474\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_\
        );

    \I__4210\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26468\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__26468\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__26465\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15_cascade_\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__26459\,
            I => \N__26456\
        );

    \I__4205\ : Span4Mux_v
    port map (
            O => \N__26456\,
            I => \N__26453\
        );

    \I__4204\ : Odrv4
    port map (
            O => \N__26453\,
            I => \phase_controller_inst2.stoper_hc.un6_running_17\
        );

    \I__4203\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26444\
        );

    \I__4202\ : InMux
    port map (
            O => \N__26449\,
            I => \N__26444\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__26444\,
            I => \elapsed_time_ns_1_RNIQ3ND11_0_22\
        );

    \I__4200\ : CascadeMux
    port map (
            O => \N__26441\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_\
        );

    \I__4199\ : InMux
    port map (
            O => \N__26438\,
            I => \N__26432\
        );

    \I__4198\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26432\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__26432\,
            I => \elapsed_time_ns_1_RNIR4ND11_0_23\
        );

    \I__4196\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26426\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__26426\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__26423\,
            I => \elapsed_time_ns_1_RNIL13KD1_0_9_cascade_\
        );

    \I__4193\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__26417\,
            I => \elapsed_time_ns_1_RNI1BND11_0_29\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__26414\,
            I => \elapsed_time_ns_1_RNI1BND11_0_29_cascade_\
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__26411\,
            I => \N__26408\
        );

    \I__4189\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26405\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__26405\,
            I => \elapsed_time_ns_1_RNIT6ND11_0_25\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26396\
        );

    \I__4186\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26396\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__26396\,
            I => \elapsed_time_ns_1_RNI0AND11_0_28\
        );

    \I__4184\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26389\
        );

    \I__4183\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26386\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__26389\,
            I => \elapsed_time_ns_1_RNIV8ND11_0_27\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__26386\,
            I => \elapsed_time_ns_1_RNIV8ND11_0_27\
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__26381\,
            I => \elapsed_time_ns_1_RNIT6ND11_0_25_cascade_\
        );

    \I__4179\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26374\
        );

    \I__4178\ : InMux
    port map (
            O => \N__26377\,
            I => \N__26371\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__26374\,
            I => \elapsed_time_ns_1_RNIU7ND11_0_26\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__26371\,
            I => \elapsed_time_ns_1_RNIU7ND11_0_26\
        );

    \I__4175\ : InMux
    port map (
            O => \N__26366\,
            I => \N__26360\
        );

    \I__4174\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26352\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26352\
        );

    \I__4172\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26352\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__26360\,
            I => \N__26349\
        );

    \I__4170\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26346\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__26352\,
            I => \N__26343\
        );

    \I__4168\ : Span4Mux_v
    port map (
            O => \N__26349\,
            I => \N__26340\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26337\
        );

    \I__4166\ : Span4Mux_h
    port map (
            O => \N__26343\,
            I => \N__26334\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__26340\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4164\ : Odrv12
    port map (
            O => \N__26337\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4163\ : Odrv4
    port map (
            O => \N__26334\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__26327\,
            I => \N__26324\
        );

    \I__4161\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26321\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__26321\,
            I => \N__26318\
        );

    \I__4159\ : Odrv4
    port map (
            O => \N__26318\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__4157\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26309\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__26309\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__26306\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc5_cascade_\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__26303\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26295\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26299\,
            I => \N__26292\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26289\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__26295\,
            I => \N__26286\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__26292\,
            I => \N__26283\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__26289\,
            I => \N__26280\
        );

    \I__4147\ : Span4Mux_h
    port map (
            O => \N__26286\,
            I => \N__26275\
        );

    \I__4146\ : Span4Mux_h
    port map (
            O => \N__26283\,
            I => \N__26270\
        );

    \I__4145\ : Span4Mux_h
    port map (
            O => \N__26280\,
            I => \N__26270\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26265\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26265\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__26275\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__26270\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__26265\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4139\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26255\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__26252\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__26249\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23_cascade_\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__26246\,
            I => \N__26243\
        );

    \I__4134\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26240\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__26240\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__26237\,
            I => \N__26233\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26236\,
            I => \N__26230\
        );

    \I__4130\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26227\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__26230\,
            I => \N__26222\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__26227\,
            I => \N__26219\
        );

    \I__4127\ : InMux
    port map (
            O => \N__26226\,
            I => \N__26216\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26225\,
            I => \N__26212\
        );

    \I__4125\ : Span4Mux_h
    port map (
            O => \N__26222\,
            I => \N__26207\
        );

    \I__4124\ : Span4Mux_h
    port map (
            O => \N__26219\,
            I => \N__26207\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26216\,
            I => \N__26204\
        );

    \I__4122\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26201\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__26212\,
            I => \N__26198\
        );

    \I__4120\ : Odrv4
    port map (
            O => \N__26207\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__26204\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__26201\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4117\ : Odrv4
    port map (
            O => \N__26198\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__26189\,
            I => \N__26186\
        );

    \I__4115\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26183\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__26183\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__26180\,
            I => \N__26177\
        );

    \I__4112\ : InMux
    port map (
            O => \N__26177\,
            I => \N__26172\
        );

    \I__4111\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26169\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26166\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__26172\,
            I => \N__26162\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__26169\,
            I => \N__26159\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__26166\,
            I => \N__26156\
        );

    \I__4106\ : InMux
    port map (
            O => \N__26165\,
            I => \N__26153\
        );

    \I__4105\ : Span4Mux_h
    port map (
            O => \N__26162\,
            I => \N__26150\
        );

    \I__4104\ : Span4Mux_v
    port map (
            O => \N__26159\,
            I => \N__26145\
        );

    \I__4103\ : Span4Mux_v
    port map (
            O => \N__26156\,
            I => \N__26145\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26153\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4101\ : Odrv4
    port map (
            O => \N__26150\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4100\ : Odrv4
    port map (
            O => \N__26145\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4099\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26135\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__26135\,
            I => \N__26132\
        );

    \I__4097\ : Span4Mux_h
    port map (
            O => \N__26132\,
            I => \N__26129\
        );

    \I__4096\ : Odrv4
    port map (
            O => \N__26129\,
            I => \current_shift_inst.PI_CTRL.integrator_i_2\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__26126\,
            I => \N__26122\
        );

    \I__4094\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26118\
        );

    \I__4093\ : InMux
    port map (
            O => \N__26122\,
            I => \N__26115\
        );

    \I__4092\ : InMux
    port map (
            O => \N__26121\,
            I => \N__26112\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__26118\,
            I => \N__26109\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__26115\,
            I => \N__26106\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__26112\,
            I => \N__26103\
        );

    \I__4088\ : Span4Mux_h
    port map (
            O => \N__26109\,
            I => \N__26096\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__26106\,
            I => \N__26096\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__26103\,
            I => \N__26093\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26088\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26088\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__26096\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__26093\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__26088\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__26081\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_\
        );

    \I__4079\ : InMux
    port map (
            O => \N__26078\,
            I => \N__26075\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__26075\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__26072\,
            I => \N__26068\
        );

    \I__4076\ : InMux
    port map (
            O => \N__26071\,
            I => \N__26065\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26062\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__26065\,
            I => \N__26058\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26062\,
            I => \N__26055\
        );

    \I__4072\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26050\
        );

    \I__4071\ : Span4Mux_v
    port map (
            O => \N__26058\,
            I => \N__26045\
        );

    \I__4070\ : Span4Mux_v
    port map (
            O => \N__26055\,
            I => \N__26045\
        );

    \I__4069\ : InMux
    port map (
            O => \N__26054\,
            I => \N__26042\
        );

    \I__4068\ : InMux
    port map (
            O => \N__26053\,
            I => \N__26039\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__26050\,
            I => \N__26036\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__26045\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__26042\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__26039\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__26036\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__26027\,
            I => \N__26024\
        );

    \I__4061\ : InMux
    port map (
            O => \N__26024\,
            I => \N__26021\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__26021\,
            I => \N__26018\
        );

    \I__4059\ : Odrv4
    port map (
            O => \N__26018\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__26015\,
            I => \N__26010\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__26014\,
            I => \N__26007\
        );

    \I__4056\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26002\
        );

    \I__4055\ : InMux
    port map (
            O => \N__26010\,
            I => \N__25999\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26007\,
            I => \N__25994\
        );

    \I__4053\ : InMux
    port map (
            O => \N__26006\,
            I => \N__25994\
        );

    \I__4052\ : InMux
    port map (
            O => \N__26005\,
            I => \N__25991\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__26002\,
            I => \N__25988\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__25999\,
            I => \N__25985\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__25994\,
            I => \N__25980\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25980\
        );

    \I__4047\ : Span4Mux_h
    port map (
            O => \N__25988\,
            I => \N__25973\
        );

    \I__4046\ : Span4Mux_h
    port map (
            O => \N__25985\,
            I => \N__25973\
        );

    \I__4045\ : Span4Mux_v
    port map (
            O => \N__25980\,
            I => \N__25973\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__25973\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__25970\,
            I => \N__25967\
        );

    \I__4042\ : InMux
    port map (
            O => \N__25967\,
            I => \N__25964\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__25964\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__25961\,
            I => \N__25958\
        );

    \I__4039\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25955\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__25955\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\
        );

    \I__4037\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25949\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__25949\,
            I => \N__25945\
        );

    \I__4035\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25942\
        );

    \I__4034\ : Span4Mux_h
    port map (
            O => \N__25945\,
            I => \N__25937\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__25942\,
            I => \N__25937\
        );

    \I__4032\ : Span4Mux_h
    port map (
            O => \N__25937\,
            I => \N__25931\
        );

    \I__4031\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25928\
        );

    \I__4030\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25923\
        );

    \I__4029\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25923\
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__25931\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__25928\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__25923\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__4024\ : InMux
    port map (
            O => \N__25913\,
            I => \N__25910\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__25910\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__25907\,
            I => \N__25903\
        );

    \I__4021\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25900\
        );

    \I__4020\ : InMux
    port map (
            O => \N__25903\,
            I => \N__25897\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__25900\,
            I => \N__25894\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__25897\,
            I => \N__25891\
        );

    \I__4017\ : Span4Mux_h
    port map (
            O => \N__25894\,
            I => \N__25883\
        );

    \I__4016\ : Span4Mux_h
    port map (
            O => \N__25891\,
            I => \N__25883\
        );

    \I__4015\ : InMux
    port map (
            O => \N__25890\,
            I => \N__25880\
        );

    \I__4014\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25877\
        );

    \I__4013\ : InMux
    port map (
            O => \N__25888\,
            I => \N__25874\
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__25883\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__25880\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__25877\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__25874\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__25865\,
            I => \N__25862\
        );

    \I__4007\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25859\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__25859\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\
        );

    \I__4005\ : InMux
    port map (
            O => \N__25856\,
            I => \N__25852\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25855\,
            I => \N__25849\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__25852\,
            I => \N__25846\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__25849\,
            I => \N__25843\
        );

    \I__4001\ : Span4Mux_h
    port map (
            O => \N__25846\,
            I => \N__25835\
        );

    \I__4000\ : Span4Mux_h
    port map (
            O => \N__25843\,
            I => \N__25835\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25832\
        );

    \I__3998\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25829\
        );

    \I__3997\ : InMux
    port map (
            O => \N__25840\,
            I => \N__25826\
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__25835\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__25832\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__25829\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__25826\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__25817\,
            I => \N__25814\
        );

    \I__3991\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25811\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__25808\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__25805\,
            I => \N__25802\
        );

    \I__3987\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25799\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__25799\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\
        );

    \I__3985\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25792\
        );

    \I__3984\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25789\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__25792\,
            I => \N__25786\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__25789\,
            I => \N__25782\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__25786\,
            I => \N__25779\
        );

    \I__3980\ : InMux
    port map (
            O => \N__25785\,
            I => \N__25776\
        );

    \I__3979\ : Span4Mux_h
    port map (
            O => \N__25782\,
            I => \N__25769\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__25779\,
            I => \N__25769\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__25776\,
            I => \N__25766\
        );

    \I__3976\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25761\
        );

    \I__3975\ : InMux
    port map (
            O => \N__25774\,
            I => \N__25761\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__25769\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__25766\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__25761\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3971\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__25751\,
            I => \N__25747\
        );

    \I__3969\ : InMux
    port map (
            O => \N__25750\,
            I => \N__25743\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__25747\,
            I => \N__25740\
        );

    \I__3967\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25737\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__25743\,
            I => \N__25732\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__25740\,
            I => \N__25727\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__25737\,
            I => \N__25727\
        );

    \I__3963\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25722\
        );

    \I__3962\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25722\
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__25732\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__25727\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__25722\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__25715\,
            I => \N__25710\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__25714\,
            I => \N__25707\
        );

    \I__3956\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25704\
        );

    \I__3955\ : InMux
    port map (
            O => \N__25710\,
            I => \N__25701\
        );

    \I__3954\ : InMux
    port map (
            O => \N__25707\,
            I => \N__25698\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__25704\,
            I => \N__25694\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__25701\,
            I => \N__25691\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__25698\,
            I => \N__25688\
        );

    \I__3950\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25684\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__25694\,
            I => \N__25681\
        );

    \I__3948\ : Span4Mux_v
    port map (
            O => \N__25691\,
            I => \N__25676\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__25688\,
            I => \N__25676\
        );

    \I__3946\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25673\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__25684\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__25681\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__25676\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__25673\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3941\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25661\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__25661\,
            I => \N__25658\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__25658\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\
        );

    \I__3938\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25651\
        );

    \I__3937\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25648\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__25651\,
            I => \N__25645\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__25648\,
            I => \N__25642\
        );

    \I__3934\ : Span4Mux_v
    port map (
            O => \N__25645\,
            I => \N__25639\
        );

    \I__3933\ : Span4Mux_h
    port map (
            O => \N__25642\,
            I => \N__25636\
        );

    \I__3932\ : Span4Mux_h
    port map (
            O => \N__25639\,
            I => \N__25633\
        );

    \I__3931\ : Odrv4
    port map (
            O => \N__25636\,
            I => \current_shift_inst.PI_CTRL.N_72\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__25633\,
            I => \current_shift_inst.PI_CTRL.N_72\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__25628\,
            I => \N__25625\
        );

    \I__3928\ : InMux
    port map (
            O => \N__25625\,
            I => \N__25622\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__25622\,
            I => \N__25619\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__25619\,
            I => \current_shift_inst.PI_CTRL.integrator_i_25\
        );

    \I__3925\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25612\
        );

    \I__3924\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25609\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__25612\,
            I => \N__25606\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__25609\,
            I => \N__25603\
        );

    \I__3921\ : Span4Mux_v
    port map (
            O => \N__25606\,
            I => \N__25600\
        );

    \I__3920\ : Span4Mux_h
    port map (
            O => \N__25603\,
            I => \N__25597\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__25600\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__25597\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__3916\ : InMux
    port map (
            O => \N__25589\,
            I => \N__25586\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__25586\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__25583\,
            I => \N__25580\
        );

    \I__3913\ : InMux
    port map (
            O => \N__25580\,
            I => \N__25577\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__25577\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__25574\,
            I => \N__25571\
        );

    \I__3910\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25568\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__25568\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__25565\,
            I => \N__25562\
        );

    \I__3907\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25559\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__25559\,
            I => \N__25555\
        );

    \I__3905\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25552\
        );

    \I__3904\ : Span4Mux_h
    port map (
            O => \N__25555\,
            I => \N__25549\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__25552\,
            I => \N__25541\
        );

    \I__3902\ : Span4Mux_h
    port map (
            O => \N__25549\,
            I => \N__25541\
        );

    \I__3901\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25536\
        );

    \I__3900\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25536\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25546\,
            I => \N__25533\
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__25541\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__25536\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__25533\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__25526\,
            I => \N__25523\
        );

    \I__3894\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__25520\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\
        );

    \I__3892\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25514\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__25514\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__25511\,
            I => \N__25506\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__25510\,
            I => \N__25502\
        );

    \I__3888\ : InMux
    port map (
            O => \N__25509\,
            I => \N__25497\
        );

    \I__3887\ : InMux
    port map (
            O => \N__25506\,
            I => \N__25497\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25505\,
            I => \N__25494\
        );

    \I__3885\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25491\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__25497\,
            I => \N__25486\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__25494\,
            I => \N__25481\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__25491\,
            I => \N__25481\
        );

    \I__3881\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25476\
        );

    \I__3880\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25476\
        );

    \I__3879\ : Odrv4
    port map (
            O => \N__25486\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3878\ : Odrv12
    port map (
            O => \N__25481\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__25476\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__25469\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__3874\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25460\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__25460\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__25457\,
            I => \N__25454\
        );

    \I__3871\ : InMux
    port map (
            O => \N__25454\,
            I => \N__25451\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__25451\,
            I => \N__25448\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__25448\,
            I => \current_shift_inst.PI_CTRL.integrator_i_4\
        );

    \I__3868\ : InMux
    port map (
            O => \N__25445\,
            I => \N__25442\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__25442\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__25439\,
            I => \N__25436\
        );

    \I__3865\ : InMux
    port map (
            O => \N__25436\,
            I => \N__25433\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__25433\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__3863\ : InMux
    port map (
            O => \N__25430\,
            I => \N__25427\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__25427\,
            I => \N__25424\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__25424\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__3860\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25418\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__25418\,
            I => \N__25415\
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__25415\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__3857\ : InMux
    port map (
            O => \N__25412\,
            I => \N__25409\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__25409\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__25406\,
            I => \N__25403\
        );

    \I__3854\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__25400\,
            I => \N__25397\
        );

    \I__3852\ : Odrv12
    port map (
            O => \N__25397\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__3850\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25388\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__3848\ : Odrv4
    port map (
            O => \N__25385\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\
        );

    \I__3847\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25375\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__25381\,
            I => \N__25372\
        );

    \I__3845\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25367\
        );

    \I__3844\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25367\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25378\,
            I => \N__25364\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25375\,
            I => \N__25361\
        );

    \I__3841\ : InMux
    port map (
            O => \N__25372\,
            I => \N__25358\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__25367\,
            I => \N__25355\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__25364\,
            I => \N__25352\
        );

    \I__3838\ : Span4Mux_v
    port map (
            O => \N__25361\,
            I => \N__25349\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__25358\,
            I => \N__25346\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__25355\,
            I => \N__25341\
        );

    \I__3835\ : Span4Mux_h
    port map (
            O => \N__25352\,
            I => \N__25341\
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__25349\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__25346\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__25341\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__25334\,
            I => \N__25331\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25328\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\
        );

    \I__3828\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25321\
        );

    \I__3827\ : InMux
    port map (
            O => \N__25324\,
            I => \N__25318\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__25321\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__25318\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25310\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__25310\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__3822\ : InMux
    port map (
            O => \N__25307\,
            I => \N__25304\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__25304\,
            I => \N__25301\
        );

    \I__3820\ : Odrv4
    port map (
            O => \N__25301\,
            I => \phase_controller_inst2.stoper_hc.un6_running_16\
        );

    \I__3819\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25294\
        );

    \I__3818\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25291\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__25294\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25291\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__25286\,
            I => \N__25283\
        );

    \I__3814\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25280\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__25280\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25273\
        );

    \I__3811\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25270\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__25273\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__25270\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__25265\,
            I => \N__25262\
        );

    \I__3807\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25259\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__25259\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\
        );

    \I__3805\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25253\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__25253\,
            I => \N__25250\
        );

    \I__3803\ : Span4Mux_v
    port map (
            O => \N__25250\,
            I => \N__25247\
        );

    \I__3802\ : Odrv4
    port map (
            O => \N__25247\,
            I => \phase_controller_inst2.stoper_hc.un6_running_18\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25244\,
            I => \N__25240\
        );

    \I__3800\ : InMux
    port map (
            O => \N__25243\,
            I => \N__25237\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__25240\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__25237\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__25232\,
            I => \N__25229\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25226\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__25226\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25223\,
            I => \N__25219\
        );

    \I__3793\ : InMux
    port map (
            O => \N__25222\,
            I => \N__25216\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__25219\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__25216\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3790\ : CascadeMux
    port map (
            O => \N__25211\,
            I => \N__25208\
        );

    \I__3789\ : InMux
    port map (
            O => \N__25208\,
            I => \N__25205\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__25205\,
            I => \N__25202\
        );

    \I__3787\ : Odrv12
    port map (
            O => \N__25202\,
            I => \phase_controller_inst2.stoper_hc.un6_running_19\
        );

    \I__3786\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25196\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__25196\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\
        );

    \I__3784\ : InMux
    port map (
            O => \N__25193\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_19\
        );

    \I__3783\ : IoInMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__25187\,
            I => \N__25184\
        );

    \I__3781\ : Span12Mux_s1_v
    port map (
            O => \N__25184\,
            I => \N__25181\
        );

    \I__3780\ : Odrv12
    port map (
            O => \N__25181\,
            I => s3_phy_c
        );

    \I__3779\ : InMux
    port map (
            O => \N__25178\,
            I => \N__25175\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__25175\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\
        );

    \I__3777\ : CascadeMux
    port map (
            O => \N__25172\,
            I => \N__25169\
        );

    \I__3776\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25166\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__25166\,
            I => \N__25163\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__25163\,
            I => \phase_controller_inst2.stoper_hc.un6_running_8\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25156\
        );

    \I__3772\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25153\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__25156\,
            I => \N__25150\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__25153\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__25150\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3768\ : InMux
    port map (
            O => \N__25145\,
            I => \N__25142\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__25142\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__3766\ : CascadeMux
    port map (
            O => \N__25139\,
            I => \N__25136\
        );

    \I__3765\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25133\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__25133\,
            I => \N__25130\
        );

    \I__3763\ : Odrv12
    port map (
            O => \N__25130\,
            I => \phase_controller_inst2.stoper_hc.un6_running_9\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25127\,
            I => \N__25123\
        );

    \I__3761\ : InMux
    port map (
            O => \N__25126\,
            I => \N__25120\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__25123\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__25120\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25115\,
            I => \N__25112\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__25112\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__3756\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25106\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__25106\,
            I => \N__25103\
        );

    \I__3754\ : Odrv12
    port map (
            O => \N__25103\,
            I => \phase_controller_inst2.stoper_hc.un6_running_10\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25096\
        );

    \I__3752\ : InMux
    port map (
            O => \N__25099\,
            I => \N__25093\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__25096\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__25093\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__25088\,
            I => \N__25085\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25085\,
            I => \N__25082\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__25082\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__3746\ : InMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__3744\ : Span4Mux_v
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__25070\,
            I => \phase_controller_inst2.stoper_hc.un6_running_11\
        );

    \I__3742\ : InMux
    port map (
            O => \N__25067\,
            I => \N__25063\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25060\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__25063\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__25060\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__3737\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__25049\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__25046\,
            I => \N__25043\
        );

    \I__3734\ : InMux
    port map (
            O => \N__25043\,
            I => \N__25040\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__25040\,
            I => \N__25037\
        );

    \I__3732\ : Odrv12
    port map (
            O => \N__25037\,
            I => \phase_controller_inst2.stoper_hc.un6_running_12\
        );

    \I__3731\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25030\
        );

    \I__3730\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25027\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__25030\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__25027\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3727\ : InMux
    port map (
            O => \N__25022\,
            I => \N__25019\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__25019\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__3725\ : InMux
    port map (
            O => \N__25016\,
            I => \N__25013\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__25013\,
            I => \N__25010\
        );

    \I__3723\ : Odrv12
    port map (
            O => \N__25010\,
            I => \phase_controller_inst2.stoper_hc.un6_running_13\
        );

    \I__3722\ : InMux
    port map (
            O => \N__25007\,
            I => \N__25003\
        );

    \I__3721\ : InMux
    port map (
            O => \N__25006\,
            I => \N__25000\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25003\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__25000\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__24995\,
            I => \N__24992\
        );

    \I__3717\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__24989\,
            I => \N__24986\
        );

    \I__3715\ : Odrv4
    port map (
            O => \N__24986\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__3714\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24980\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__24980\,
            I => \N__24977\
        );

    \I__3712\ : Odrv12
    port map (
            O => \N__24977\,
            I => \phase_controller_inst2.stoper_hc.un6_running_14\
        );

    \I__3711\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24970\
        );

    \I__3710\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24967\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__24970\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__24967\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3707\ : CascadeMux
    port map (
            O => \N__24962\,
            I => \N__24959\
        );

    \I__3706\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24956\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__24956\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__24953\,
            I => \N__24946\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__24952\,
            I => \N__24935\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__24951\,
            I => \N__24932\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__24950\,
            I => \N__24929\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__24949\,
            I => \N__24926\
        );

    \I__3699\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24922\
        );

    \I__3698\ : InMux
    port map (
            O => \N__24945\,
            I => \N__24919\
        );

    \I__3697\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24910\
        );

    \I__3696\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24910\
        );

    \I__3695\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24910\
        );

    \I__3694\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24910\
        );

    \I__3693\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24897\
        );

    \I__3692\ : InMux
    port map (
            O => \N__24939\,
            I => \N__24897\
        );

    \I__3691\ : InMux
    port map (
            O => \N__24938\,
            I => \N__24897\
        );

    \I__3690\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24897\
        );

    \I__3689\ : InMux
    port map (
            O => \N__24932\,
            I => \N__24897\
        );

    \I__3688\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24897\
        );

    \I__3687\ : InMux
    port map (
            O => \N__24926\,
            I => \N__24892\
        );

    \I__3686\ : InMux
    port map (
            O => \N__24925\,
            I => \N__24892\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__24922\,
            I => \N__24889\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__24919\,
            I => \N__24886\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__24910\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__24897\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__24892\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__24889\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__3679\ : Odrv12
    port map (
            O => \N__24886\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__3677\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24856\
        );

    \I__3676\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24856\
        );

    \I__3675\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24853\
        );

    \I__3674\ : InMux
    port map (
            O => \N__24869\,
            I => \N__24846\
        );

    \I__3673\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24846\
        );

    \I__3672\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24846\
        );

    \I__3671\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24839\
        );

    \I__3670\ : InMux
    port map (
            O => \N__24865\,
            I => \N__24839\
        );

    \I__3669\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24839\
        );

    \I__3668\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24836\
        );

    \I__3667\ : InMux
    port map (
            O => \N__24862\,
            I => \N__24831\
        );

    \I__3666\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24831\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__24856\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__24853\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__24846\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__24839\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__24836\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__24831\,
            I => \phase_controller_inst1.stoper_hc.N_327\
        );

    \I__3659\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24815\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24812\
        );

    \I__3657\ : Span4Mux_v
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__24809\,
            I => \phase_controller_inst2.stoper_hc.un6_running_1\
        );

    \I__3655\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24802\
        );

    \I__3654\ : CascadeMux
    port map (
            O => \N__24805\,
            I => \N__24798\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__24802\,
            I => \N__24795\
        );

    \I__3652\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24792\
        );

    \I__3651\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24789\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__24795\,
            I => \N__24786\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__24792\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__24789\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__24786\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__24779\,
            I => \N__24776\
        );

    \I__3645\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__24773\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__3643\ : InMux
    port map (
            O => \N__24770\,
            I => \N__24767\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__24767\,
            I => \phase_controller_inst2.stoper_hc.un6_running_2\
        );

    \I__3641\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24760\
        );

    \I__3640\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24757\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__24760\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__24757\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3637\ : CascadeMux
    port map (
            O => \N__24752\,
            I => \N__24749\
        );

    \I__3636\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24746\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__24746\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__3634\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24739\
        );

    \I__3633\ : InMux
    port map (
            O => \N__24742\,
            I => \N__24736\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__24739\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__24736\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3630\ : InMux
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__24728\,
            I => \N__24725\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__24725\,
            I => \N__24722\
        );

    \I__3627\ : Odrv4
    port map (
            O => \N__24722\,
            I => \phase_controller_inst2.stoper_hc.un6_running_3\
        );

    \I__3626\ : CascadeMux
    port map (
            O => \N__24719\,
            I => \N__24716\
        );

    \I__3625\ : InMux
    port map (
            O => \N__24716\,
            I => \N__24713\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__24713\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__3623\ : InMux
    port map (
            O => \N__24710\,
            I => \N__24707\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__24707\,
            I => \N__24703\
        );

    \I__3621\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24700\
        );

    \I__3620\ : Sp12to4
    port map (
            O => \N__24703\,
            I => \N__24697\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__24700\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3618\ : Odrv12
    port map (
            O => \N__24697\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3617\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24689\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__24689\,
            I => \phase_controller_inst2.stoper_hc.un6_running_4\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__24686\,
            I => \N__24683\
        );

    \I__3614\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24680\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__24680\,
            I => \N__24677\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__24677\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__3611\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24671\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__3609\ : Odrv4
    port map (
            O => \N__24668\,
            I => \phase_controller_inst2.stoper_hc.un6_running_5\
        );

    \I__3608\ : InMux
    port map (
            O => \N__24665\,
            I => \N__24661\
        );

    \I__3607\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24658\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__24661\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__24658\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3604\ : CascadeMux
    port map (
            O => \N__24653\,
            I => \N__24650\
        );

    \I__3603\ : InMux
    port map (
            O => \N__24650\,
            I => \N__24647\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__24647\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__3601\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24640\
        );

    \I__3600\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24637\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__24640\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__24637\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__24632\,
            I => \N__24629\
        );

    \I__3596\ : InMux
    port map (
            O => \N__24629\,
            I => \N__24626\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__24626\,
            I => \N__24623\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__24623\,
            I => \phase_controller_inst2.stoper_hc.un6_running_6\
        );

    \I__3593\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__24617\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__24614\,
            I => \N__24611\
        );

    \I__3590\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__24605\,
            I => \phase_controller_inst2.stoper_hc.un6_running_7\
        );

    \I__3587\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24598\
        );

    \I__3586\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24595\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__24598\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__24595\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3583\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24587\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__24587\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__24584\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_\
        );

    \I__3580\ : CascadeMux
    port map (
            O => \N__24581\,
            I => \N__24577\
        );

    \I__3579\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24573\
        );

    \I__3578\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24570\
        );

    \I__3577\ : InMux
    port map (
            O => \N__24576\,
            I => \N__24567\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__24573\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__24570\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__24567\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__24560\,
            I => \elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_\
        );

    \I__3572\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24552\
        );

    \I__3571\ : InMux
    port map (
            O => \N__24556\,
            I => \N__24547\
        );

    \I__3570\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24547\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__24552\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__24547\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__24542\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__24539\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6_cascade_\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__24536\,
            I => \N__24532\
        );

    \I__3564\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24529\
        );

    \I__3563\ : InMux
    port map (
            O => \N__24532\,
            I => \N__24526\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__24529\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__24526\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__24521\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\
        );

    \I__3559\ : InMux
    port map (
            O => \N__24518\,
            I => \N__24512\
        );

    \I__3558\ : InMux
    port map (
            O => \N__24517\,
            I => \N__24509\
        );

    \I__3557\ : InMux
    port map (
            O => \N__24516\,
            I => \N__24504\
        );

    \I__3556\ : InMux
    port map (
            O => \N__24515\,
            I => \N__24504\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__24512\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__24509\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__24504\,
            I => \elapsed_time_ns_1_RNIDP2KD1_0_1\
        );

    \I__3552\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24493\
        );

    \I__3551\ : InMux
    port map (
            O => \N__24496\,
            I => \N__24490\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__24493\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__24490\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__24485\,
            I => \elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_\
        );

    \I__3547\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__24479\,
            I => \N__24476\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__24476\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__24473\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9_cascade_\
        );

    \I__3543\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24462\
        );

    \I__3542\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24462\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__24468\,
            I => \N__24454\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__24467\,
            I => \N__24451\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__24462\,
            I => \N__24446\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24441\
        );

    \I__3537\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24441\
        );

    \I__3536\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24438\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24458\,
            I => \N__24431\
        );

    \I__3534\ : InMux
    port map (
            O => \N__24457\,
            I => \N__24431\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24431\
        );

    \I__3532\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24428\
        );

    \I__3531\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24423\
        );

    \I__3530\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24423\
        );

    \I__3529\ : Sp12to4
    port map (
            O => \N__24446\,
            I => \N__24418\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__24441\,
            I => \N__24418\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__24438\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__24431\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__24428\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__24423\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__3523\ : Odrv12
    port map (
            O => \N__24418\,
            I => \phase_controller_inst1.stoper_hc.N_315\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__24407\,
            I => \N__24403\
        );

    \I__3521\ : InMux
    port map (
            O => \N__24406\,
            I => \N__24400\
        );

    \I__3520\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24397\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__24400\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__24397\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__24392\,
            I => \phase_controller_inst1.stoper_hc.N_283_cascade_\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24385\
        );

    \I__3515\ : InMux
    port map (
            O => \N__24388\,
            I => \N__24382\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__24385\,
            I => \phase_controller_inst1.stoper_hc.N_307\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__24382\,
            I => \phase_controller_inst1.stoper_hc.N_307\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24374\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24374\,
            I => \N__24371\
        );

    \I__3510\ : Span4Mux_h
    port map (
            O => \N__24371\,
            I => \N__24368\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__24368\,
            I => \phase_controller_inst1.stoper_hc.un6_running_7\
        );

    \I__3508\ : CEMux
    port map (
            O => \N__24365\,
            I => \N__24357\
        );

    \I__3507\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24343\
        );

    \I__3506\ : InMux
    port map (
            O => \N__24363\,
            I => \N__24343\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24343\
        );

    \I__3504\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24343\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24360\,
            I => \N__24340\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24357\,
            I => \N__24337\
        );

    \I__3501\ : CEMux
    port map (
            O => \N__24356\,
            I => \N__24333\
        );

    \I__3500\ : InMux
    port map (
            O => \N__24355\,
            I => \N__24314\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24354\,
            I => \N__24314\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24314\
        );

    \I__3497\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24314\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__24343\,
            I => \N__24309\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__24340\,
            I => \N__24309\
        );

    \I__3494\ : Span4Mux_v
    port map (
            O => \N__24337\,
            I => \N__24306\
        );

    \I__3493\ : CEMux
    port map (
            O => \N__24336\,
            I => \N__24303\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24300\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24293\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24331\,
            I => \N__24293\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24293\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24284\
        );

    \I__3487\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24284\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24284\
        );

    \I__3485\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24284\
        );

    \I__3484\ : InMux
    port map (
            O => \N__24325\,
            I => \N__24277\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24277\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24323\,
            I => \N__24277\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24270\
        );

    \I__3480\ : Span4Mux_v
    port map (
            O => \N__24309\,
            I => \N__24270\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__24306\,
            I => \N__24270\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__24303\,
            I => \N__24263\
        );

    \I__3477\ : Span4Mux_v
    port map (
            O => \N__24300\,
            I => \N__24263\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__24293\,
            I => \N__24263\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__24284\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__24277\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__3473\ : Odrv4
    port map (
            O => \N__24270\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__24263\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__24254\,
            I => \elapsed_time_ns_1_RNI62CED1_0_19_cascade_\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__24251\,
            I => \phase_controller_inst1.stoper_hc.N_315_cascade_\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__24248\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_\
        );

    \I__3468\ : InMux
    port map (
            O => \N__24245\,
            I => \N__24242\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__24242\,
            I => \N__24239\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__24239\,
            I => \phase_controller_inst1.stoper_hc.un6_running_9\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__24236\,
            I => \N__24233\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24230\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24227\
        );

    \I__3462\ : Odrv12
    port map (
            O => \N__24227\,
            I => \phase_controller_inst1.stoper_hc.un6_running_13\
        );

    \I__3461\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24221\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24221\,
            I => \N__24218\
        );

    \I__3459\ : Span4Mux_h
    port map (
            O => \N__24218\,
            I => \N__24215\
        );

    \I__3458\ : Odrv4
    port map (
            O => \N__24215\,
            I => \phase_controller_inst1.stoper_hc.un6_running_19\
        );

    \I__3457\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24209\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__3455\ : Span4Mux_h
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__24203\,
            I => \phase_controller_inst1.stoper_hc.un6_running_18\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24197\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__3451\ : Span4Mux_v
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__24191\,
            I => \phase_controller_inst1.stoper_hc.un6_running_17\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24185\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__24185\,
            I => \N__24182\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__24182\,
            I => \phase_controller_inst1.stoper_hc.un6_running_16\
        );

    \I__3446\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24176\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24173\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__24173\,
            I => \phase_controller_inst1.stoper_hc.un6_running_15\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__24170\,
            I => \N__24167\
        );

    \I__3442\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24164\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__24164\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__3440\ : InMux
    port map (
            O => \N__24161\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\
        );

    \I__3439\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24155\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__24155\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__3437\ : InMux
    port map (
            O => \N__24152\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24149\,
            I => \bfn_9_12_0_\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24146\,
            I => \N__24143\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__24143\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__24140\,
            I => \N__24137\
        );

    \I__3432\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24130\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24136\,
            I => \N__24130\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24127\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__24130\,
            I => \N__24123\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N__24120\
        );

    \I__3427\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24117\
        );

    \I__3426\ : Span4Mux_v
    port map (
            O => \N__24123\,
            I => \N__24114\
        );

    \I__3425\ : Odrv12
    port map (
            O => \N__24120\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24117\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__24114\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__24107\,
            I => \N__24104\
        );

    \I__3421\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24101\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__24101\,
            I => \current_shift_inst.PI_CTRL.integrator_i_29\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__24098\,
            I => \N__24093\
        );

    \I__3418\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24088\
        );

    \I__3417\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24088\
        );

    \I__3416\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24085\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__24088\,
            I => \N__24081\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24085\,
            I => \N__24078\
        );

    \I__3413\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24075\
        );

    \I__3412\ : Span4Mux_h
    port map (
            O => \N__24081\,
            I => \N__24072\
        );

    \I__3411\ : Odrv12
    port map (
            O => \N__24078\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__24075\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3409\ : Odrv4
    port map (
            O => \N__24072\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24065\,
            I => \N__24062\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__24062\,
            I => \current_shift_inst.PI_CTRL.integrator_i_28\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__24059\,
            I => \N__24056\
        );

    \I__3405\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24053\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__24053\,
            I => \N__24050\
        );

    \I__3403\ : Odrv4
    port map (
            O => \N__24050\,
            I => \current_shift_inst.PI_CTRL.integrator_i_15\
        );

    \I__3402\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24042\
        );

    \I__3401\ : InMux
    port map (
            O => \N__24046\,
            I => \N__24035\
        );

    \I__3400\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24035\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__24042\,
            I => \N__24032\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__24041\,
            I => \N__24029\
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__24040\,
            I => \N__24026\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__24035\,
            I => \N__24023\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__24032\,
            I => \N__24020\
        );

    \I__3394\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24017\
        );

    \I__3393\ : InMux
    port map (
            O => \N__24026\,
            I => \N__24014\
        );

    \I__3392\ : Span4Mux_v
    port map (
            O => \N__24023\,
            I => \N__24011\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__24020\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__24017\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__24014\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__24011\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3387\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23999\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__23999\,
            I => \N__23996\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__23996\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\
        );

    \I__3384\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23990\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__23990\,
            I => \N__23987\
        );

    \I__3382\ : Span4Mux_h
    port map (
            O => \N__23987\,
            I => \N__23984\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__23984\,
            I => \current_shift_inst.PI_CTRL.integrator_i_22\
        );

    \I__3380\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__23978\,
            I => \N__23975\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__23975\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__3377\ : InMux
    port map (
            O => \N__23972\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__23969\,
            I => \N__23966\
        );

    \I__3375\ : InMux
    port map (
            O => \N__23966\,
            I => \N__23963\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__23963\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__3373\ : InMux
    port map (
            O => \N__23960\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\
        );

    \I__3372\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23954\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__23954\,
            I => \N__23951\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__23948\,
            I => \current_shift_inst.PI_CTRL.integrator_i_23\
        );

    \I__3368\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23942\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__23942\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__3366\ : InMux
    port map (
            O => \N__23939\,
            I => \bfn_9_11_0_\
        );

    \I__3365\ : InMux
    port map (
            O => \N__23936\,
            I => \N__23933\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__23933\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__3363\ : InMux
    port map (
            O => \N__23930\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__3361\ : InMux
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__23921\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__3359\ : InMux
    port map (
            O => \N__23918\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__23915\,
            I => \N__23912\
        );

    \I__3357\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23909\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__23909\,
            I => \N__23906\
        );

    \I__3355\ : Odrv12
    port map (
            O => \N__23906\,
            I => \current_shift_inst.PI_CTRL.integrator_i_26\
        );

    \I__3354\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23900\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__23900\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__3352\ : InMux
    port map (
            O => \N__23897\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\
        );

    \I__3351\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23891\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__23891\,
            I => \N__23888\
        );

    \I__3349\ : Span4Mux_h
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__23885\,
            I => \current_shift_inst.PI_CTRL.integrator_i_27\
        );

    \I__3347\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23876\
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__23876\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__3344\ : InMux
    port map (
            O => \N__23873\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\
        );

    \I__3343\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23867\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__23867\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__3341\ : InMux
    port map (
            O => \N__23864\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23861\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\
        );

    \I__3339\ : InMux
    port map (
            O => \N__23858\,
            I => \N__23855\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__23855\,
            I => \N__23852\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__23852\,
            I => \current_shift_inst.PI_CTRL.integrator_i_14\
        );

    \I__3336\ : InMux
    port map (
            O => \N__23849\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\
        );

    \I__3335\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__23843\,
            I => \N__23840\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__23840\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__3332\ : InMux
    port map (
            O => \N__23837\,
            I => \bfn_9_10_0_\
        );

    \I__3331\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23831\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__23831\,
            I => \N__23828\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__23828\,
            I => \current_shift_inst.PI_CTRL.integrator_i_16\
        );

    \I__3328\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23822\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__23822\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__3326\ : InMux
    port map (
            O => \N__23819\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\
        );

    \I__3325\ : InMux
    port map (
            O => \N__23816\,
            I => \N__23813\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__23813\,
            I => \N__23810\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__23810\,
            I => \current_shift_inst.PI_CTRL.integrator_i_17\
        );

    \I__3322\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23804\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__23804\,
            I => \N__23801\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__23801\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__3319\ : InMux
    port map (
            O => \N__23798\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\
        );

    \I__3318\ : InMux
    port map (
            O => \N__23795\,
            I => \N__23792\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__23792\,
            I => \N__23789\
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__23789\,
            I => \current_shift_inst.PI_CTRL.integrator_i_18\
        );

    \I__3315\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23783\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__23783\,
            I => \N__23780\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__23780\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__3312\ : InMux
    port map (
            O => \N__23777\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\
        );

    \I__3311\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23771\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__23771\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__3309\ : InMux
    port map (
            O => \N__23768\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\
        );

    \I__3308\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23762\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__23762\,
            I => \N__23759\
        );

    \I__3306\ : Odrv12
    port map (
            O => \N__23759\,
            I => \current_shift_inst.PI_CTRL.integrator_i_20\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__3304\ : InMux
    port map (
            O => \N__23753\,
            I => \N__23750\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__23750\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__3302\ : InMux
    port map (
            O => \N__23747\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\
        );

    \I__3301\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23741\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__23741\,
            I => \current_shift_inst.PI_CTRL.integrator_i_5\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__23738\,
            I => \N__23735\
        );

    \I__3298\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23732\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__23732\,
            I => \N__23729\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__23729\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__23726\,
            I => \N__23723\
        );

    \I__3294\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23720\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__23720\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__3292\ : InMux
    port map (
            O => \N__23717\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\
        );

    \I__3291\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23711\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__23711\,
            I => \N__23708\
        );

    \I__3289\ : Span4Mux_v
    port map (
            O => \N__23708\,
            I => \N__23705\
        );

    \I__3288\ : Odrv4
    port map (
            O => \N__23705\,
            I => \current_shift_inst.PI_CTRL.integrator_i_6\
        );

    \I__3287\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23699\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__23699\,
            I => \N__23696\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__23696\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__3284\ : InMux
    port map (
            O => \N__23693\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\
        );

    \I__3283\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23687\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__23687\,
            I => \current_shift_inst.PI_CTRL.integrator_i_7\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__23684\,
            I => \N__23681\
        );

    \I__3280\ : InMux
    port map (
            O => \N__23681\,
            I => \N__23678\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__23678\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\
        );

    \I__3278\ : InMux
    port map (
            O => \N__23675\,
            I => \N__23672\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__23672\,
            I => \N__23669\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__23669\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3275\ : InMux
    port map (
            O => \N__23666\,
            I => \bfn_9_9_0_\
        );

    \I__3274\ : InMux
    port map (
            O => \N__23663\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\
        );

    \I__3273\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23657\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23654\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__23651\,
            I => \current_shift_inst.PI_CTRL.integrator_i_9\
        );

    \I__3269\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23645\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__23642\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__3266\ : InMux
    port map (
            O => \N__23639\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__3263\ : Span4Mux_h
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__23627\,
            I => \current_shift_inst.PI_CTRL.integrator_i_10\
        );

    \I__3261\ : InMux
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__23618\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__3258\ : InMux
    port map (
            O => \N__23615\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\
        );

    \I__3257\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__23609\,
            I => \current_shift_inst.PI_CTRL.integrator_i_11\
        );

    \I__3255\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__23603\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__3253\ : InMux
    port map (
            O => \N__23600\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23597\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\
        );

    \I__3251\ : IoInMux
    port map (
            O => \N__23594\,
            I => \N__23591\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__23591\,
            I => \N__23588\
        );

    \I__3249\ : Span4Mux_s2_v
    port map (
            O => \N__23588\,
            I => \N__23585\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__23582\,
            I => \delay_measurement_inst.delay_tr_timer.N_434_i\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__23573\,
            I => \N__23568\
        );

    \I__3243\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23565\
        );

    \I__3242\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23562\
        );

    \I__3241\ : Span4Mux_v
    port map (
            O => \N__23568\,
            I => \N__23557\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__23565\,
            I => \N__23557\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__23562\,
            I => \N__23554\
        );

    \I__3238\ : Span4Mux_h
    port map (
            O => \N__23557\,
            I => \N__23551\
        );

    \I__3237\ : Span4Mux_h
    port map (
            O => \N__23554\,
            I => \N__23548\
        );

    \I__3236\ : Span4Mux_v
    port map (
            O => \N__23551\,
            I => \N__23545\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__23548\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__23545\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3233\ : InMux
    port map (
            O => \N__23540\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\
        );

    \I__3232\ : InMux
    port map (
            O => \N__23537\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\
        );

    \I__3231\ : InMux
    port map (
            O => \N__23534\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\
        );

    \I__3230\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23528\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__23528\,
            I => \current_shift_inst.PI_CTRL.integrator_i_3\
        );

    \I__3228\ : InMux
    port map (
            O => \N__23525\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\
        );

    \I__3227\ : InMux
    port map (
            O => \N__23522\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\
        );

    \I__3226\ : InMux
    port map (
            O => \N__23519\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__3225\ : InMux
    port map (
            O => \N__23516\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__3224\ : InMux
    port map (
            O => \N__23513\,
            I => \bfn_8_21_0_\
        );

    \I__3223\ : InMux
    port map (
            O => \N__23510\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__3222\ : InMux
    port map (
            O => \N__23507\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__3221\ : InMux
    port map (
            O => \N__23504\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__3220\ : InMux
    port map (
            O => \N__23501\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__3219\ : InMux
    port map (
            O => \N__23498\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__3218\ : InMux
    port map (
            O => \N__23495\,
            I => \bfn_8_20_0_\
        );

    \I__3217\ : InMux
    port map (
            O => \N__23492\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__3216\ : InMux
    port map (
            O => \N__23489\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__3215\ : InMux
    port map (
            O => \N__23486\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__3214\ : InMux
    port map (
            O => \N__23483\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__3213\ : InMux
    port map (
            O => \N__23480\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__3212\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23474\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__3210\ : Span4Mux_v
    port map (
            O => \N__23471\,
            I => \N__23468\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__23468\,
            I => \phase_controller_inst1.stoper_hc.un6_running_5\
        );

    \I__3208\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23462\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__23462\,
            I => \N__23459\
        );

    \I__3206\ : Span4Mux_v
    port map (
            O => \N__23459\,
            I => \N__23456\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__23456\,
            I => \phase_controller_inst1.stoper_hc.un6_running_8\
        );

    \I__3204\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23450\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__3202\ : Span4Mux_v
    port map (
            O => \N__23447\,
            I => \N__23444\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__23444\,
            I => \phase_controller_inst1.stoper_hc.un6_running_3\
        );

    \I__3200\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23438\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__23438\,
            I => \N__23435\
        );

    \I__3198\ : Span4Mux_v
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__23432\,
            I => \phase_controller_inst1.stoper_hc.un6_running_1\
        );

    \I__3196\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23426\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__23426\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23423\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__23420\,
            I => \N__23417\
        );

    \I__3192\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23414\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23411\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__23411\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21\
        );

    \I__3189\ : InMux
    port map (
            O => \N__23408\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__3188\ : InMux
    port map (
            O => \N__23405\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23402\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__3186\ : InMux
    port map (
            O => \N__23399\,
            I => \N__23396\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__3184\ : Span4Mux_v
    port map (
            O => \N__23393\,
            I => \N__23390\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__23390\,
            I => \phase_controller_inst1.stoper_hc.un6_running_6\
        );

    \I__3182\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23384\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__23384\,
            I => \N__23381\
        );

    \I__3180\ : Span4Mux_v
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__23378\,
            I => \phase_controller_inst1.stoper_hc.un6_running_2\
        );

    \I__3178\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23372\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__23372\,
            I => \N__23369\
        );

    \I__3176\ : Span4Mux_v
    port map (
            O => \N__23369\,
            I => \N__23366\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__23366\,
            I => \phase_controller_inst1.stoper_hc.un6_running_4\
        );

    \I__3174\ : InMux
    port map (
            O => \N__23363\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23356\
        );

    \I__3172\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23353\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__23356\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__23353\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__23348\,
            I => \N__23344\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__23347\,
            I => \N__23340\
        );

    \I__3167\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23337\
        );

    \I__3166\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23334\
        );

    \I__3165\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23331\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__23337\,
            I => \N__23326\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__23334\,
            I => \N__23326\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__23331\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__23326\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3160\ : InMux
    port map (
            O => \N__23321\,
            I => \N__23317\
        );

    \I__3159\ : InMux
    port map (
            O => \N__23320\,
            I => \N__23314\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23317\,
            I => \phase_controller_inst1.stoper_hc.running_1_sqmuxa\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__23314\,
            I => \phase_controller_inst1.stoper_hc.running_1_sqmuxa\
        );

    \I__3156\ : InMux
    port map (
            O => \N__23309\,
            I => \N__23306\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__23303\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__3153\ : InMux
    port map (
            O => \N__23300\,
            I => \N__23296\
        );

    \I__3152\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23293\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__23296\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__23293\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO\
        );

    \I__3149\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23284\
        );

    \I__3148\ : InMux
    port map (
            O => \N__23287\,
            I => \N__23281\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__23284\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__23281\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__23276\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23270\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__23270\,
            I => \N__23267\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__23267\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTIZ0Z1\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23259\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23254\
        );

    \I__3139\ : InMux
    port map (
            O => \N__23262\,
            I => \N__23254\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__23259\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__23254\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__3136\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23243\
        );

    \I__3135\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23240\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23247\,
            I => \N__23235\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23235\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__23243\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__23240\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__23235\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23224\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23221\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__23224\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__23221\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3125\ : InMux
    port map (
            O => \N__23216\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__3124\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23209\
        );

    \I__3123\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23206\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__23209\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__23206\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23201\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23194\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23191\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__23194\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__23191\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23186\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__3114\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23179\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23176\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__23179\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__23176\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23171\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23164\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23161\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23164\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__23161\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3105\ : InMux
    port map (
            O => \N__23156\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__3104\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23149\
        );

    \I__3103\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23146\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__23149\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__23146\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3100\ : InMux
    port map (
            O => \N__23141\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__3099\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23134\
        );

    \I__3098\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23131\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__23134\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__23131\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3095\ : InMux
    port map (
            O => \N__23126\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23119\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23122\,
            I => \N__23116\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__23119\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23116\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3090\ : InMux
    port map (
            O => \N__23111\,
            I => \bfn_8_15_0_\
        );

    \I__3089\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23104\
        );

    \I__3088\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23101\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__23104\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__23101\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23096\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23089\
        );

    \I__3083\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23086\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__23089\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__23086\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23081\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__23078\,
            I => \N__23075\
        );

    \I__3078\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23071\
        );

    \I__3077\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23068\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__23071\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__23068\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3074\ : InMux
    port map (
            O => \N__23063\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23056\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23053\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__23056\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__23053\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3069\ : InMux
    port map (
            O => \N__23048\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__3068\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23041\
        );

    \I__3067\ : InMux
    port map (
            O => \N__23044\,
            I => \N__23038\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__23041\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__23038\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3064\ : InMux
    port map (
            O => \N__23033\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__3063\ : InMux
    port map (
            O => \N__23030\,
            I => \N__23026\
        );

    \I__3062\ : InMux
    port map (
            O => \N__23029\,
            I => \N__23023\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__23026\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__23023\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3059\ : InMux
    port map (
            O => \N__23018\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__3058\ : InMux
    port map (
            O => \N__23015\,
            I => \N__23011\
        );

    \I__3057\ : InMux
    port map (
            O => \N__23014\,
            I => \N__23008\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__23011\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__23008\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3054\ : InMux
    port map (
            O => \N__23003\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__3053\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22996\
        );

    \I__3052\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22993\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__22996\,
            I => \N__22988\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__22993\,
            I => \N__22988\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__22988\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3048\ : InMux
    port map (
            O => \N__22985\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22978\
        );

    \I__3046\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22975\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__22978\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__22975\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3043\ : InMux
    port map (
            O => \N__22970\,
            I => \bfn_8_14_0_\
        );

    \I__3042\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22964\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__22964\,
            I => \N__22961\
        );

    \I__3040\ : Span4Mux_h
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__22958\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__22955\,
            I => \N__22946\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__22954\,
            I => \N__22942\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__22953\,
            I => \N__22938\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__22952\,
            I => \N__22930\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__22951\,
            I => \N__22926\
        );

    \I__3033\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22908\
        );

    \I__3032\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22908\
        );

    \I__3031\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22908\
        );

    \I__3030\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22908\
        );

    \I__3029\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22908\
        );

    \I__3028\ : InMux
    port map (
            O => \N__22941\,
            I => \N__22908\
        );

    \I__3027\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22908\
        );

    \I__3026\ : InMux
    port map (
            O => \N__22937\,
            I => \N__22908\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__22936\,
            I => \N__22905\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__22935\,
            I => \N__22901\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__22934\,
            I => \N__22897\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__22933\,
            I => \N__22893\
        );

    \I__3021\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22883\
        );

    \I__3020\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22883\
        );

    \I__3019\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22883\
        );

    \I__3018\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22883\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__22908\,
            I => \N__22880\
        );

    \I__3016\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22863\
        );

    \I__3015\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22863\
        );

    \I__3014\ : InMux
    port map (
            O => \N__22901\,
            I => \N__22863\
        );

    \I__3013\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22863\
        );

    \I__3012\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22863\
        );

    \I__3011\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22863\
        );

    \I__3010\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22863\
        );

    \I__3009\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22863\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__22883\,
            I => \N__22860\
        );

    \I__3007\ : Span4Mux_v
    port map (
            O => \N__22880\,
            I => \N__22855\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__22863\,
            I => \N__22855\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__22860\,
            I => \N__22852\
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__22855\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3003\ : Odrv4
    port map (
            O => \N__22852\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3002\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22843\
        );

    \I__3001\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22840\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__22843\,
            I => \current_shift_inst.PI_CTRL.N_74_16\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__22840\,
            I => \current_shift_inst.PI_CTRL.N_74_16\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__22835\,
            I => \N__22832\
        );

    \I__2997\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22828\
        );

    \I__2996\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22825\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__22828\,
            I => \N__22822\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__22825\,
            I => \current_shift_inst.PI_CTRL.N_74_21\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__22822\,
            I => \current_shift_inst.PI_CTRL.N_74_21\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__22817\,
            I => \current_shift_inst.PI_CTRL.N_103_cascade_\
        );

    \I__2991\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22811\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__22811\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__22808\,
            I => \N__22805\
        );

    \I__2988\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22799\
        );

    \I__2987\ : InMux
    port map (
            O => \N__22804\,
            I => \N__22799\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__22799\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__22796\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__2984\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22786\
        );

    \I__2983\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22786\
        );

    \I__2982\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22783\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__22786\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__22783\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__2979\ : InMux
    port map (
            O => \N__22778\,
            I => \N__22775\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__2977\ : Odrv12
    port map (
            O => \N__22772\,
            I => il_max_comp1_c
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__2975\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22763\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__22763\,
            I => \N__22758\
        );

    \I__2973\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22753\
        );

    \I__2972\ : InMux
    port map (
            O => \N__22761\,
            I => \N__22753\
        );

    \I__2971\ : Span4Mux_h
    port map (
            O => \N__22758\,
            I => \N__22748\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__22753\,
            I => \N__22745\
        );

    \I__2969\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22740\
        );

    \I__2968\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22740\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__22748\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__22745\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__22740\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__22733\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_\
        );

    \I__2963\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__22727\,
            I => \phase_controller_inst2.start_timer_hc_RNOZ0Z_0\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__22724\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__2959\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__22715\,
            I => \N__22712\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__22712\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__22709\,
            I => \N__22706\
        );

    \I__2955\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22703\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__22703\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \N__22697\
        );

    \I__2952\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22694\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__22694\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__22691\,
            I => \N__22688\
        );

    \I__2949\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22685\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__22685\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__2946\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__22676\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__2944\ : InMux
    port map (
            O => \N__22673\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_19\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__22670\,
            I => \N__22667\
        );

    \I__2942\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__22664\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__22661\,
            I => \N__22658\
        );

    \I__2939\ : InMux
    port map (
            O => \N__22658\,
            I => \N__22655\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__22655\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__2937\ : CascadeMux
    port map (
            O => \N__22652\,
            I => \N__22649\
        );

    \I__2936\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22646\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__22646\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__2934\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22640\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__22640\,
            I => \N__22637\
        );

    \I__2932\ : Span4Mux_v
    port map (
            O => \N__22637\,
            I => \N__22634\
        );

    \I__2931\ : Odrv4
    port map (
            O => \N__22634\,
            I => \phase_controller_inst1.stoper_hc.un6_running_10\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__22631\,
            I => \N__22628\
        );

    \I__2929\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22625\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__22625\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__2927\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22619\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__22619\,
            I => \N__22616\
        );

    \I__2925\ : Span4Mux_h
    port map (
            O => \N__22616\,
            I => \N__22613\
        );

    \I__2924\ : Odrv4
    port map (
            O => \N__22613\,
            I => \phase_controller_inst1.stoper_hc.un6_running_11\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__22610\,
            I => \N__22607\
        );

    \I__2922\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22604\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__22604\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__2920\ : InMux
    port map (
            O => \N__22601\,
            I => \N__22598\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__22598\,
            I => \N__22595\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__22595\,
            I => \N__22592\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__22592\,
            I => \phase_controller_inst1.stoper_hc.un6_running_12\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__22583\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__2913\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22577\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__22577\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__2911\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22571\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__22571\,
            I => \N__22568\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__22565\,
            I => \phase_controller_inst1.stoper_hc.un6_running_14\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__2906\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22556\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__22556\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__2903\ : InMux
    port map (
            O => \N__22550\,
            I => \N__22547\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__22547\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__22544\,
            I => \N__22541\
        );

    \I__2900\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__22538\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__2897\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__22529\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__22526\,
            I => \N__22523\
        );

    \I__2894\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22520\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__22520\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__22517\,
            I => \N__22514\
        );

    \I__2891\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22511\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__22511\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__2888\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__22502\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__2886\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__22496\,
            I => \N__22493\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__22493\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__22490\,
            I => \N__22487\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22484\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22481\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__22481\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2879\ : InMux
    port map (
            O => \N__22478\,
            I => \N__22475\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__22475\,
            I => \N__22472\
        );

    \I__2877\ : Span4Mux_h
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__22469\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2875\ : InMux
    port map (
            O => \N__22466\,
            I => \N__22463\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__22463\,
            I => \N__22460\
        );

    \I__2873\ : Odrv12
    port map (
            O => \N__22460\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2872\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22454\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__22454\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\
        );

    \I__2870\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__2868\ : Span4Mux_v
    port map (
            O => \N__22445\,
            I => \N__22442\
        );

    \I__2867\ : Odrv4
    port map (
            O => \N__22442\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__22436\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\
        );

    \I__2864\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22430\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__22430\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\
        );

    \I__2862\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__22424\,
            I => \current_shift_inst.PI_CTRL.N_62\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__22421\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_\
        );

    \I__2859\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__22415\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__2857\ : InMux
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__22409\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__2854\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__2852\ : Span4Mux_v
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__2851\ : Odrv4
    port map (
            O => \N__22394\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22391\,
            I => \N__22388\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__22388\,
            I => \N__22385\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__22385\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22379\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__22379\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22373\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__22373\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__22370\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__22367\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__22364\,
            I => \current_shift_inst.PI_CTRL.N_75_cascade_\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22355\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22355\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__22355\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22352\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__2835\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22340\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22340\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__22340\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2832\ : InMux
    port map (
            O => \N__22337\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2831\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__22331\,
            I => \N__22327\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22324\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__22327\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__22324\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2826\ : InMux
    port map (
            O => \N__22319\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22307\
        );

    \I__2823\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22307\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22304\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__22304\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22301\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22295\,
            I => \N__22291\
        );

    \I__2817\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22288\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__22291\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__22288\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22283\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2813\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__22277\,
            I => \N__22273\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__22276\,
            I => \N__22270\
        );

    \I__2810\ : Span4Mux_h
    port map (
            O => \N__22273\,
            I => \N__22267\
        );

    \I__2809\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22264\
        );

    \I__2808\ : Odrv4
    port map (
            O => \N__22267\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__22264\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22259\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2805\ : InMux
    port map (
            O => \N__22256\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2804\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22249\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__22252\,
            I => \N__22245\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__22249\,
            I => \N__22236\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22227\
        );

    \I__2800\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22227\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22227\
        );

    \I__2798\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22227\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22224\
        );

    \I__2796\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22221\
        );

    \I__2795\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22216\
        );

    \I__2794\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22216\
        );

    \I__2793\ : Span4Mux_v
    port map (
            O => \N__22236\,
            I => \N__22204\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__22227\,
            I => \N__22204\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__22224\,
            I => \N__22204\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__22221\,
            I => \N__22204\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__22216\,
            I => \N__22204\
        );

    \I__2788\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22201\
        );

    \I__2787\ : Span4Mux_v
    port map (
            O => \N__22204\,
            I => \N__22196\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__22201\,
            I => \N__22196\
        );

    \I__2785\ : Span4Mux_h
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__22193\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2783\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__22181\,
            I => \il_max_comp2_D1\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22171\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22174\,
            I => \N__22168\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__22171\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__22168\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22163\,
            I => \bfn_5_11_0_\
        );

    \I__2773\ : InMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__22157\,
            I => \N__22153\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22150\
        );

    \I__2770\ : Odrv4
    port map (
            O => \N__22153\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__22150\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22145\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__22139\,
            I => \N__22135\
        );

    \I__2765\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22132\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__22135\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__22132\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2762\ : InMux
    port map (
            O => \N__22127\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22118\
        );

    \I__2760\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22118\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__22118\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2758\ : InMux
    port map (
            O => \N__22115\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__22112\,
            I => \N__22108\
        );

    \I__2756\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22103\
        );

    \I__2755\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22103\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__22103\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2753\ : InMux
    port map (
            O => \N__22100\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__22097\,
            I => \N__22093\
        );

    \I__2751\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22088\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22088\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__22088\,
            I => \N__22085\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__22085\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2747\ : InMux
    port map (
            O => \N__22082\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2746\ : InMux
    port map (
            O => \N__22079\,
            I => \N__22073\
        );

    \I__2745\ : InMux
    port map (
            O => \N__22078\,
            I => \N__22073\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__22073\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2743\ : InMux
    port map (
            O => \N__22070\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22063\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22060\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__22063\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__22060\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2738\ : InMux
    port map (
            O => \N__22055\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__2736\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__22046\,
            I => \N__22042\
        );

    \I__2734\ : InMux
    port map (
            O => \N__22045\,
            I => \N__22039\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__22042\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__22039\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2731\ : InMux
    port map (
            O => \N__22034\,
            I => \bfn_5_12_0_\
        );

    \I__2730\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22026\
        );

    \I__2729\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22023\
        );

    \I__2728\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22020\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__22026\,
            I => \N__22017\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__22023\,
            I => \N__22012\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__22020\,
            I => \N__22012\
        );

    \I__2724\ : Span4Mux_h
    port map (
            O => \N__22017\,
            I => \N__22009\
        );

    \I__2723\ : Odrv12
    port map (
            O => \N__22012\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2722\ : Odrv4
    port map (
            O => \N__22009\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2721\ : InMux
    port map (
            O => \N__22004\,
            I => \bfn_5_10_0_\
        );

    \I__2720\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__21998\,
            I => \N__21993\
        );

    \I__2718\ : InMux
    port map (
            O => \N__21997\,
            I => \N__21990\
        );

    \I__2717\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21987\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__21993\,
            I => \N__21984\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__21990\,
            I => \N__21979\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21979\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__21984\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2712\ : Odrv12
    port map (
            O => \N__21979\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2711\ : InMux
    port map (
            O => \N__21974\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2710\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21965\
        );

    \I__2709\ : InMux
    port map (
            O => \N__21970\,
            I => \N__21965\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__21965\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2707\ : InMux
    port map (
            O => \N__21962\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2706\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__21956\,
            I => \N__21952\
        );

    \I__2704\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21949\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__21952\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__21949\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2701\ : InMux
    port map (
            O => \N__21944\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__2699\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__21935\,
            I => \N__21931\
        );

    \I__2697\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21928\
        );

    \I__2696\ : Odrv4
    port map (
            O => \N__21931\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__21928\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2694\ : InMux
    port map (
            O => \N__21923\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2693\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21916\
        );

    \I__2692\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21913\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__21916\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__21913\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2689\ : InMux
    port map (
            O => \N__21908\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2688\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21901\
        );

    \I__2687\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21898\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__21901\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__21898\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2684\ : InMux
    port map (
            O => \N__21893\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2683\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21886\
        );

    \I__2682\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21883\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__21886\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__21883\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2679\ : InMux
    port map (
            O => \N__21878\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2678\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__21872\,
            I => \N__21869\
        );

    \I__2676\ : Odrv12
    port map (
            O => \N__21869\,
            I => il_max_comp2_c
        );

    \I__2675\ : InMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__21863\,
            I => \N__21860\
        );

    \I__2673\ : Odrv12
    port map (
            O => \N__21860\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2672\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__2670\ : Odrv12
    port map (
            O => \N__21851\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2669\ : InMux
    port map (
            O => \N__21848\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2668\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__21842\,
            I => \N__21839\
        );

    \I__2666\ : Odrv12
    port map (
            O => \N__21839\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2665\ : InMux
    port map (
            O => \N__21836\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2664\ : InMux
    port map (
            O => \N__21833\,
            I => \N__21828\
        );

    \I__2663\ : InMux
    port map (
            O => \N__21832\,
            I => \N__21825\
        );

    \I__2662\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21822\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__21828\,
            I => \N__21817\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__21825\,
            I => \N__21817\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__21822\,
            I => \N__21812\
        );

    \I__2658\ : Span4Mux_v
    port map (
            O => \N__21817\,
            I => \N__21812\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__21812\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2656\ : InMux
    port map (
            O => \N__21809\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2655\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21802\
        );

    \I__2654\ : InMux
    port map (
            O => \N__21805\,
            I => \N__21798\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__21802\,
            I => \N__21794\
        );

    \I__2652\ : InMux
    port map (
            O => \N__21801\,
            I => \N__21791\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__21798\,
            I => \N__21788\
        );

    \I__2650\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21785\
        );

    \I__2649\ : Span4Mux_v
    port map (
            O => \N__21794\,
            I => \N__21780\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__21791\,
            I => \N__21780\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__21788\,
            I => \N__21777\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__21785\,
            I => \N__21774\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__21780\,
            I => \N__21771\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__21777\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__21774\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__21771\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2641\ : InMux
    port map (
            O => \N__21764\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__2639\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21753\
        );

    \I__2638\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21750\
        );

    \I__2637\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21747\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__21753\,
            I => \N__21740\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__21750\,
            I => \N__21740\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__21747\,
            I => \N__21740\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__21737\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2631\ : InMux
    port map (
            O => \N__21734\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2630\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21726\
        );

    \I__2629\ : InMux
    port map (
            O => \N__21730\,
            I => \N__21723\
        );

    \I__2628\ : InMux
    port map (
            O => \N__21729\,
            I => \N__21720\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__21726\,
            I => \N__21715\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__21723\,
            I => \N__21715\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__21720\,
            I => \N__21712\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__21715\,
            I => \N__21709\
        );

    \I__2623\ : Span4Mux_h
    port map (
            O => \N__21712\,
            I => \N__21706\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__21709\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__21706\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2620\ : InMux
    port map (
            O => \N__21701\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2619\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21693\
        );

    \I__2618\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21690\
        );

    \I__2617\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21687\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__21693\,
            I => \N__21684\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__21690\,
            I => \N__21679\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__21687\,
            I => \N__21679\
        );

    \I__2613\ : Span4Mux_h
    port map (
            O => \N__21684\,
            I => \N__21676\
        );

    \I__2612\ : Span4Mux_h
    port map (
            O => \N__21679\,
            I => \N__21673\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__21676\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__21673\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2609\ : InMux
    port map (
            O => \N__21668\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2608\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__21659\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__2605\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__2603\ : Span4Mux_h
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__21647\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__2600\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21638\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21638\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__2598\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__21632\,
            I => \N__21629\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__21629\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__2595\ : InMux
    port map (
            O => \N__21626\,
            I => \N__21623\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__21623\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__2593\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21617\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__21617\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2591\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__2589\ : Span4Mux_h
    port map (
            O => \N__21608\,
            I => \N__21605\
        );

    \I__2588\ : Odrv4
    port map (
            O => \N__21605\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__2587\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21599\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__21599\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__2585\ : InMux
    port map (
            O => \N__21596\,
            I => \N__21593\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__21593\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2583\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21577\
        );

    \I__2582\ : InMux
    port map (
            O => \N__21589\,
            I => \N__21577\
        );

    \I__2581\ : InMux
    port map (
            O => \N__21588\,
            I => \N__21572\
        );

    \I__2580\ : InMux
    port map (
            O => \N__21587\,
            I => \N__21572\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21586\,
            I => \N__21561\
        );

    \I__2578\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21561\
        );

    \I__2577\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21561\
        );

    \I__2576\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21561\
        );

    \I__2575\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21561\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__21577\,
            I => \N__21558\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__21572\,
            I => \N__21555\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21551\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__21558\,
            I => \N__21546\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__21555\,
            I => \N__21546\
        );

    \I__2569\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21543\
        );

    \I__2568\ : Span4Mux_v
    port map (
            O => \N__21551\,
            I => \N__21540\
        );

    \I__2567\ : Span4Mux_v
    port map (
            O => \N__21546\,
            I => \N__21537\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__21543\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__21540\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__21537\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2563\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21522\
        );

    \I__2562\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21522\
        );

    \I__2561\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21517\
        );

    \I__2560\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21517\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__21522\,
            I => \N__21509\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__21517\,
            I => \N__21506\
        );

    \I__2557\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21495\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21495\
        );

    \I__2555\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21495\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21495\
        );

    \I__2553\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21495\
        );

    \I__2552\ : Span4Mux_v
    port map (
            O => \N__21509\,
            I => \N__21490\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__21506\,
            I => \N__21490\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__21495\,
            I => \N__21487\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__21490\,
            I => \N__21483\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__21487\,
            I => \N__21480\
        );

    \I__2547\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21477\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__21483\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__21480\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__21477\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \N__21465\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__21469\,
            I => \N__21461\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__21468\,
            I => \N__21458\
        );

    \I__2540\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21453\
        );

    \I__2539\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21453\
        );

    \I__2538\ : InMux
    port map (
            O => \N__21461\,
            I => \N__21448\
        );

    \I__2537\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21448\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__21453\,
            I => \N__21445\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__21448\,
            I => \N__21442\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__21445\,
            I => \N__21431\
        );

    \I__2533\ : Span4Mux_h
    port map (
            O => \N__21442\,
            I => \N__21428\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21423\
        );

    \I__2531\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21423\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__21439\,
            I => \N__21420\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__21438\,
            I => \N__21417\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__21437\,
            I => \N__21414\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__21436\,
            I => \N__21411\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__21435\,
            I => \N__21408\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__21434\,
            I => \N__21405\
        );

    \I__2524\ : Span4Mux_h
    port map (
            O => \N__21431\,
            I => \N__21398\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__21428\,
            I => \N__21398\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__21423\,
            I => \N__21398\
        );

    \I__2521\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21392\
        );

    \I__2520\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21385\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21385\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21385\
        );

    \I__2517\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21380\
        );

    \I__2516\ : InMux
    port map (
            O => \N__21405\,
            I => \N__21380\
        );

    \I__2515\ : Span4Mux_v
    port map (
            O => \N__21398\,
            I => \N__21376\
        );

    \I__2514\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21369\
        );

    \I__2513\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21369\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21369\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21362\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__21385\,
            I => \N__21362\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21362\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__21379\,
            I => \N__21359\
        );

    \I__2507\ : Span4Mux_s1_h
    port map (
            O => \N__21376\,
            I => \N__21338\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__21369\,
            I => \N__21338\
        );

    \I__2505\ : Span12Mux_v
    port map (
            O => \N__21362\,
            I => \N__21335\
        );

    \I__2504\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21332\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21329\
        );

    \I__2502\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21312\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21312\
        );

    \I__2500\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21312\
        );

    \I__2499\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21312\
        );

    \I__2498\ : InMux
    port map (
            O => \N__21353\,
            I => \N__21312\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21312\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21312\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21312\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21297\
        );

    \I__2493\ : InMux
    port map (
            O => \N__21348\,
            I => \N__21297\
        );

    \I__2492\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21297\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21297\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21345\,
            I => \N__21297\
        );

    \I__2489\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21297\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21297\
        );

    \I__2487\ : Span4Mux_v
    port map (
            O => \N__21338\,
            I => \N__21294\
        );

    \I__2486\ : Odrv12
    port map (
            O => \N__21335\,
            I => \N_19_1\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N_19_1\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__21329\,
            I => \N_19_1\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__21312\,
            I => \N_19_1\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N_19_1\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__21294\,
            I => \N_19_1\
        );

    \I__2480\ : InMux
    port map (
            O => \N__21281\,
            I => \N__21278\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21278\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__2478\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21272\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__21272\,
            I => \N__21269\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__21269\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__21260\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21254\,
            I => \N__21250\
        );

    \I__2470\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21247\
        );

    \I__2469\ : Span4Mux_h
    port map (
            O => \N__21250\,
            I => \N__21241\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__21247\,
            I => \N__21241\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21238\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__21241\,
            I => \N__21235\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__21238\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__21235\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__21230\,
            I => \N__21227\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21224\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__2460\ : Span4Mux_h
    port map (
            O => \N__21221\,
            I => \N__21217\
        );

    \I__2459\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21214\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__21217\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__21214\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__21209\,
            I => \N__21205\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__21208\,
            I => \N__21198\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21194\
        );

    \I__2453\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21191\
        );

    \I__2452\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21186\
        );

    \I__2451\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21186\
        );

    \I__2450\ : InMux
    port map (
            O => \N__21201\,
            I => \N__21183\
        );

    \I__2449\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21180\
        );

    \I__2448\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21177\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__21194\,
            I => \N__21173\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__21191\,
            I => \N__21170\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21164\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__21183\,
            I => \N__21157\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__21180\,
            I => \N__21157\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__21177\,
            I => \N__21157\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21154\
        );

    \I__2440\ : Span4Mux_v
    port map (
            O => \N__21173\,
            I => \N__21151\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__21170\,
            I => \N__21148\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21145\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21142\
        );

    \I__2436\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21139\
        );

    \I__2435\ : Span4Mux_s2_h
    port map (
            O => \N__21164\,
            I => \N__21132\
        );

    \I__2434\ : Span4Mux_h
    port map (
            O => \N__21157\,
            I => \N__21132\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__21154\,
            I => \N__21132\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__21151\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__21148\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__21145\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__21142\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__21139\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__21132\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2426\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__21116\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__2424\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21108\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21112\,
            I => \N__21105\
        );

    \I__2422\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21102\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__21108\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__21105\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__21102\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2418\ : InMux
    port map (
            O => \N__21095\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__2417\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21087\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21084\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21081\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__21087\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__21084\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__21081\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2411\ : InMux
    port map (
            O => \N__21074\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21066\
        );

    \I__2409\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21063\
        );

    \I__2408\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21060\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__21066\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__21063\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__21060\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21053\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__2403\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21045\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21049\,
            I => \N__21042\
        );

    \I__2401\ : InMux
    port map (
            O => \N__21048\,
            I => \N__21039\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__21045\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__21042\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__21039\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2397\ : InMux
    port map (
            O => \N__21032\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__2396\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21024\
        );

    \I__2395\ : InMux
    port map (
            O => \N__21028\,
            I => \N__21021\
        );

    \I__2394\ : InMux
    port map (
            O => \N__21027\,
            I => \N__21018\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__21024\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__21021\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__21018\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21011\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21008\,
            I => \N__21003\
        );

    \I__2388\ : InMux
    port map (
            O => \N__21007\,
            I => \N__21000\
        );

    \I__2387\ : InMux
    port map (
            O => \N__21006\,
            I => \N__20997\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__21003\,
            I => \N__20994\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__21000\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__20997\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__20994\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2382\ : InMux
    port map (
            O => \N__20987\,
            I => \bfn_4_14_0_\
        );

    \I__2381\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20970\
        );

    \I__2380\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20970\
        );

    \I__2379\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20970\
        );

    \I__2378\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20970\
        );

    \I__2377\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20961\
        );

    \I__2376\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20961\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__20970\,
            I => \N__20958\
        );

    \I__2374\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20949\
        );

    \I__2373\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20949\
        );

    \I__2372\ : InMux
    port map (
            O => \N__20967\,
            I => \N__20949\
        );

    \I__2371\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20949\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__20961\,
            I => \N__20946\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__20958\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__20949\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__20946\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2366\ : InMux
    port map (
            O => \N__20939\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__2365\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20931\
        );

    \I__2364\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20928\
        );

    \I__2363\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20925\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__20931\,
            I => \N__20922\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__20928\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__20925\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__20922\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__20915\,
            I => \N__20912\
        );

    \I__2357\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__20906\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__2354\ : InMux
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__20900\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2352\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__20894\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__20891\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__20888\,
            I => \pwm_generator_inst.un1_counterlto9_2_cascade_\
        );

    \I__2348\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20882\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__20882\,
            I => \pwm_generator_inst.un1_counterlt9\
        );

    \I__2346\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20874\
        );

    \I__2345\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20871\
        );

    \I__2344\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20868\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__20874\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__20871\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__20868\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2340\ : InMux
    port map (
            O => \N__20861\,
            I => \bfn_4_13_0_\
        );

    \I__2339\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20853\
        );

    \I__2338\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20850\
        );

    \I__2337\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20847\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__20853\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__20850\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__20847\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2333\ : InMux
    port map (
            O => \N__20840\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__2332\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20832\
        );

    \I__2331\ : InMux
    port map (
            O => \N__20836\,
            I => \N__20829\
        );

    \I__2330\ : InMux
    port map (
            O => \N__20835\,
            I => \N__20826\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__20832\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__20829\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__20826\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2326\ : InMux
    port map (
            O => \N__20819\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__20816\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__20810\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2322\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__20804\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2320\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20798\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__20798\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__20795\,
            I => \N__20792\
        );

    \I__2317\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20789\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__20789\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__20786\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__2314\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__20780\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2312\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__20774\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9\
        );

    \I__2310\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20768\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__20768\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2308\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20762\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__20762\,
            I => \N__20759\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__20759\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__2305\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__20753\,
            I => \N__20750\
        );

    \I__2303\ : Span12Mux_s9_v
    port map (
            O => \N__20750\,
            I => \N__20747\
        );

    \I__2302\ : Odrv12
    port map (
            O => \N__20747\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__2301\ : InMux
    port map (
            O => \N__20744\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__2300\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20738\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__20738\,
            I => \N__20735\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__20735\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__2297\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20729\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__20729\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__2295\ : InMux
    port map (
            O => \N__20726\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__2294\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20720\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__20717\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__2291\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__20711\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__2289\ : InMux
    port map (
            O => \N__20708\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__2288\ : InMux
    port map (
            O => \N__20705\,
            I => \bfn_3_18_0_\
        );

    \I__2287\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__20699\,
            I => \N__20696\
        );

    \I__2285\ : Span4Mux_v
    port map (
            O => \N__20696\,
            I => \N__20693\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__20693\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__2283\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20687\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__20687\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2281\ : InMux
    port map (
            O => \N__20684\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__2280\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20678\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__20675\,
            I => \N__20671\
        );

    \I__2277\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20668\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__20671\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__20668\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__20663\,
            I => \N__20659\
        );

    \I__2273\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20655\
        );

    \I__2272\ : InMux
    port map (
            O => \N__20659\,
            I => \N__20652\
        );

    \I__2271\ : InMux
    port map (
            O => \N__20658\,
            I => \N__20649\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__20655\,
            I => \N__20644\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__20652\,
            I => \N__20644\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__20649\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__20644\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2266\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20636\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__20636\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__2264\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__20630\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__2262\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20624\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__20624\,
            I => \N__20621\
        );

    \I__2260\ : Glb2LocalMux
    port map (
            O => \N__20621\,
            I => \N__20618\
        );

    \I__2259\ : GlobalMux
    port map (
            O => \N__20618\,
            I => clk_12mhz
        );

    \I__2258\ : IoInMux
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__2256\ : Span4Mux_s0_v
    port map (
            O => \N__20609\,
            I => \N__20606\
        );

    \I__2255\ : Sp12to4
    port map (
            O => \N__20606\,
            I => \N__20603\
        );

    \I__2254\ : Odrv12
    port map (
            O => \N__20603\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2253\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20597\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__20597\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2251\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__20591\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__2249\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20585\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__2247\ : Odrv12
    port map (
            O => \N__20582\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__2246\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20576\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__20576\,
            I => \N__20573\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__20573\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__2243\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20567\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__20567\,
            I => \N__20564\
        );

    \I__2241\ : Odrv12
    port map (
            O => \N__20564\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2240\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__20558\,
            I => \N__20555\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__20555\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__2237\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__20549\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__2235\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20543\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__20543\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__2233\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20537\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__20537\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__2231\ : InMux
    port map (
            O => \N__20534\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20528\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20525\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__20525\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__2227\ : InMux
    port map (
            O => \N__20522\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20519\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__2225\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20513\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__20513\,
            I => \N__20510\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__20510\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__2222\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20504\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__20504\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__2220\ : InMux
    port map (
            O => \N__20501\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__2219\ : CascadeMux
    port map (
            O => \N__20498\,
            I => \N__20495\
        );

    \I__2218\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20492\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__20492\,
            I => \N__20489\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__20489\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__2215\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20483\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__20483\,
            I => \N__20480\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__20480\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__2212\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20473\
        );

    \I__2211\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20470\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__20473\,
            I => \N__20467\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20464\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__20467\,
            I => \N__20461\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__20464\,
            I => \N__20458\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__20461\,
            I => \pwm_generator_inst.O_10\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__20458\,
            I => \pwm_generator_inst.O_10\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20450\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__20450\,
            I => \N__20446\
        );

    \I__2202\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20442\
        );

    \I__2201\ : Span4Mux_h
    port map (
            O => \N__20446\,
            I => \N__20439\
        );

    \I__2200\ : InMux
    port map (
            O => \N__20445\,
            I => \N__20436\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__20442\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__20439\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__20436\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__2195\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__20423\,
            I => \N__20420\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__20420\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__2192\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__20411\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__20402\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__20396\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__20387\,
            I => \N__20384\
        );

    \I__2181\ : Span4Mux_h
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__20381\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__20375\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20366\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__20366\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__2173\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__20357\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__20348\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__2167\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__20339\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2165\ : InMux
    port map (
            O => \N__20336\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2164\ : IoInMux
    port map (
            O => \N__20333\,
            I => \N__20330\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__20330\,
            I => \N__20327\
        );

    \I__2162\ : Span4Mux_s2_v
    port map (
            O => \N__20327\,
            I => \N__20324\
        );

    \I__2161\ : Sp12to4
    port map (
            O => \N__20324\,
            I => \N__20321\
        );

    \I__2160\ : Span12Mux_s10_h
    port map (
            O => \N__20321\,
            I => \N__20318\
        );

    \I__2159\ : Span12Mux_h
    port map (
            O => \N__20318\,
            I => \N__20315\
        );

    \I__2158\ : Odrv12
    port map (
            O => \N__20315\,
            I => pwm_output_c
        );

    \I__2157\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20309\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__20309\,
            I => \N__20306\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__20306\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__2154\ : InMux
    port map (
            O => \N__20303\,
            I => \N__20300\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__2152\ : Odrv4
    port map (
            O => \N__20297\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__2151\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20291\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__20291\,
            I => \N__20287\
        );

    \I__2149\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20283\
        );

    \I__2148\ : Span4Mux_h
    port map (
            O => \N__20287\,
            I => \N__20280\
        );

    \I__2147\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20277\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__20283\,
            I => pwm_duty_input_5
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__20280\,
            I => pwm_duty_input_5
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__20277\,
            I => pwm_duty_input_5
        );

    \I__2143\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20267\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__20267\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__20264\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__20261\,
            I => \N__20254\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20250\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20239\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20239\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20239\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20254\,
            I => \N__20239\
        );

    \I__2134\ : InMux
    port map (
            O => \N__20253\,
            I => \N__20239\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__20250\,
            I => \N__20236\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__20239\,
            I => \N__20228\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__20236\,
            I => \N__20228\
        );

    \I__2130\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20225\
        );

    \I__2129\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20220\
        );

    \I__2128\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20220\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__20228\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__20225\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20220\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2124\ : InMux
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__20210\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__20207\,
            I => \N__20201\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__20206\,
            I => \N__20198\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__20205\,
            I => \N__20195\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__20204\,
            I => \N__20192\
        );

    \I__2118\ : InMux
    port map (
            O => \N__20201\,
            I => \N__20179\
        );

    \I__2117\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20179\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20179\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20179\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20179\
        );

    \I__2113\ : InMux
    port map (
            O => \N__20190\,
            I => \N__20176\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__20179\,
            I => \N__20173\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__20176\,
            I => \N__20169\
        );

    \I__2110\ : Span4Mux_s3_h
    port map (
            O => \N__20173\,
            I => \N__20166\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20172\,
            I => \N__20163\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__20169\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__20166\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__20163\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__20150\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__2101\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20141\,
            I => \N__20138\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__20138\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2098\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20132\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__20132\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20123\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2093\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20116\
        );

    \I__2092\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20113\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__20116\,
            I => \N__20110\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__20113\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__20110\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__20099\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__2085\ : InMux
    port map (
            O => \N__20096\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__2084\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20089\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20086\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__20089\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__20086\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2080\ : InMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20078\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20075\,
            I => \bfn_2_18_0_\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20068\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20065\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20068\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__20065\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2073\ : InMux
    port map (
            O => \N__20060\,
            I => \N__20057\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__20057\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20054\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__2070\ : InMux
    port map (
            O => \N__20051\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__2069\ : InMux
    port map (
            O => \N__20048\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__2068\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__20042\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__2066\ : InMux
    port map (
            O => \N__20039\,
            I => \N__20036\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__20033\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2063\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__20027\,
            I => \N__20022\
        );

    \I__2061\ : InMux
    port map (
            O => \N__20026\,
            I => \N__20019\
        );

    \I__2060\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20016\
        );

    \I__2059\ : Span4Mux_h
    port map (
            O => \N__20022\,
            I => \N__20013\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__20019\,
            I => \N__20010\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__20016\,
            I => \N__20007\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__20013\,
            I => pwm_duty_input_8
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__20010\,
            I => pwm_duty_input_8
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__20007\,
            I => pwm_duty_input_8
        );

    \I__2053\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19995\
        );

    \I__2052\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19992\
        );

    \I__2051\ : InMux
    port map (
            O => \N__19998\,
            I => \N__19989\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__19995\,
            I => \N__19986\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__19992\,
            I => \N__19983\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__19989\,
            I => \N__19980\
        );

    \I__2047\ : Span4Mux_h
    port map (
            O => \N__19986\,
            I => \N__19977\
        );

    \I__2046\ : Span4Mux_h
    port map (
            O => \N__19983\,
            I => \N__19974\
        );

    \I__2045\ : Span4Mux_s1_h
    port map (
            O => \N__19980\,
            I => \N__19971\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__19977\,
            I => pwm_duty_input_9
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__19974\,
            I => pwm_duty_input_9
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__19971\,
            I => pwm_duty_input_9
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \N__19960\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__19963\,
            I => \N__19957\
        );

    \I__2039\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19953\
        );

    \I__2038\ : InMux
    port map (
            O => \N__19957\,
            I => \N__19950\
        );

    \I__2037\ : InMux
    port map (
            O => \N__19956\,
            I => \N__19947\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__19953\,
            I => \N__19942\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__19950\,
            I => \N__19942\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__19947\,
            I => \N__19939\
        );

    \I__2033\ : Span4Mux_v
    port map (
            O => \N__19942\,
            I => \N__19936\
        );

    \I__2032\ : Span4Mux_s1_h
    port map (
            O => \N__19939\,
            I => \N__19933\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__19936\,
            I => pwm_duty_input_6
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__19933\,
            I => pwm_duty_input_6
        );

    \I__2029\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__19925\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__2027\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19918\
        );

    \I__2026\ : InMux
    port map (
            O => \N__19921\,
            I => \N__19914\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__19918\,
            I => \N__19911\
        );

    \I__2024\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19908\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__19914\,
            I => \N__19905\
        );

    \I__2022\ : Span4Mux_h
    port map (
            O => \N__19911\,
            I => \N__19900\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__19908\,
            I => \N__19900\
        );

    \I__2020\ : Odrv12
    port map (
            O => \N__19905\,
            I => pwm_duty_input_7
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__19900\,
            I => pwm_duty_input_7
        );

    \I__2018\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__2016\ : Span4Mux_h
    port map (
            O => \N__19889\,
            I => \N__19886\
        );

    \I__2015\ : Span4Mux_v
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__19883\,
            I => \pwm_generator_inst.O_7\
        );

    \I__2013\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__19877\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__2011\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__2009\ : Span4Mux_h
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__2008\ : Span4Mux_v
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__19862\,
            I => \pwm_generator_inst.O_8\
        );

    \I__2006\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__19856\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__2004\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__2002\ : Span4Mux_h
    port map (
            O => \N__19847\,
            I => \N__19844\
        );

    \I__2001\ : Span4Mux_v
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__19841\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1999\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__19835\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__1997\ : InMux
    port map (
            O => \N__19832\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__1996\ : InMux
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__1994\ : Span4Mux_v
    port map (
            O => \N__19823\,
            I => \N__19819\
        );

    \I__1993\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19816\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__19819\,
            I => \N__19813\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__19816\,
            I => \N__19810\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__19813\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__19810\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1988\ : InMux
    port map (
            O => \N__19805\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__1987\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19797\
        );

    \I__1986\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19794\
        );

    \I__1985\ : InMux
    port map (
            O => \N__19800\,
            I => \N__19791\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__19797\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__19794\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__19791\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__1981\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__19778\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__1978\ : InMux
    port map (
            O => \N__19775\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__1977\ : InMux
    port map (
            O => \N__19772\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__1976\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19765\
        );

    \I__1975\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19762\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__19765\,
            I => \N__19759\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__19762\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__19759\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1971\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__1969\ : Span4Mux_h
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__19745\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__1967\ : InMux
    port map (
            O => \N__19742\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__1966\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19733\
        );

    \I__1965\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19733\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__19733\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__19730\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_\
        );

    \I__1962\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__1960\ : Span4Mux_h
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__19715\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1957\ : InMux
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__19709\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__1955\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__19700\,
            I => \N__19697\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__19694\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1950\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__19688\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__1948\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__1945\ : Span4Mux_v
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__19673\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1943\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__19667\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__1941\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__19652\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1936\ : InMux
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__19646\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__1934\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__1931\ : Span4Mux_v
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__19631\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1929\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__19625\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__1927\ : InMux
    port map (
            O => \N__19622\,
            I => \N__19619\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__19610\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1922\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__19604\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__1920\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__1918\ : Span12Mux_h
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__19592\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1916\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__19586\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__19583\,
            I => \N__19580\
        );

    \I__1913\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__19577\,
            I => \N__19574\
        );

    \I__1911\ : Span12Mux_v
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__1910\ : Odrv12
    port map (
            O => \N__19571\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1909\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__19562\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__1906\ : InMux
    port map (
            O => \N__19559\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1905\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__1902\ : Span4Mux_v
    port map (
            O => \N__19547\,
            I => \N__19544\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__19544\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1900\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19532\
        );

    \I__1899\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19529\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__19539\,
            I => \N__19526\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__19538\,
            I => \N__19522\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__19537\,
            I => \N__19519\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__19536\,
            I => \N__19516\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__19535\,
            I => \N__19513\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__19532\,
            I => \N__19510\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__19529\,
            I => \N__19507\
        );

    \I__1891\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19498\
        );

    \I__1890\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19498\
        );

    \I__1889\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19498\
        );

    \I__1888\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19498\
        );

    \I__1887\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19493\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19493\
        );

    \I__1885\ : Span4Mux_v
    port map (
            O => \N__19510\,
            I => \N__19490\
        );

    \I__1884\ : Span4Mux_h
    port map (
            O => \N__19507\,
            I => \N__19487\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__19498\,
            I => \N__19482\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__19493\,
            I => \N__19482\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__19490\,
            I => \N__19479\
        );

    \I__1880\ : Span4Mux_v
    port map (
            O => \N__19487\,
            I => \N__19476\
        );

    \I__1879\ : Span4Mux_h
    port map (
            O => \N__19482\,
            I => \N__19473\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__19479\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__19476\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__19473\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__19466\,
            I => \N__19463\
        );

    \I__1874\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__19457\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__1871\ : InMux
    port map (
            O => \N__19454\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1870\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19448\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__19448\,
            I => \N__19445\
        );

    \I__1868\ : Span4Mux_h
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__1867\ : Odrv4
    port map (
            O => \N__19442\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__1866\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19436\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__19436\,
            I => \N__19433\
        );

    \I__1864\ : Span12Mux_v
    port map (
            O => \N__19433\,
            I => \N__19430\
        );

    \I__1863\ : Odrv12
    port map (
            O => \N__19430\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1862\ : InMux
    port map (
            O => \N__19427\,
            I => \bfn_2_15_0_\
        );

    \I__1861\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19420\
        );

    \I__1860\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19417\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__19420\,
            I => \N__19414\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__19417\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__19414\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__19409\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\
        );

    \I__1855\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19400\
        );

    \I__1854\ : InMux
    port map (
            O => \N__19405\,
            I => \N__19400\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__19400\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__19397\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19391\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__19391\,
            I => \N__19388\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__19385\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__1846\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__1844\ : Span12Mux_v
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1843\ : Odrv12
    port map (
            O => \N__19370\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1842\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__19361\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19358\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1838\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__19343\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__1832\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__1830\ : Span4Mux_h
    port map (
            O => \N__19331\,
            I => \N__19328\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__19328\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__1827\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__19316\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__1824\ : InMux
    port map (
            O => \N__19313\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1823\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19307\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__19307\,
            I => \N__19304\
        );

    \I__1821\ : Span12Mux_h
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__1820\ : Odrv12
    port map (
            O => \N__19301\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__1816\ : Span4Mux_h
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__19286\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1814\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19280\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__19280\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__1812\ : InMux
    port map (
            O => \N__19277\,
            I => \bfn_2_14_0_\
        );

    \I__1811\ : InMux
    port map (
            O => \N__19274\,
            I => \N__19271\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__1809\ : Span4Mux_v
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__19262\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__1803\ : Span4Mux_h
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__19247\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19241\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__19241\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__1799\ : InMux
    port map (
            O => \N__19238\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1798\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__1796\ : Span4Mux_v
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__1795\ : Span4Mux_v
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__19223\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1793\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__19217\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19214\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__19208\,
            I => \N__19205\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__19199\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1785\ : InMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__19193\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19190\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1782\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__19175\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1777\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19169\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__19166\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__1774\ : InMux
    port map (
            O => \N__19163\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__1770\ : Span4Mux_v
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__19148\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__19145\,
            I => \N__19142\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__19136\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__1764\ : InMux
    port map (
            O => \N__19133\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__19130\,
            I => \N__19125\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19129\,
            I => \N__19116\
        );

    \I__1761\ : InMux
    port map (
            O => \N__19128\,
            I => \N__19116\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19116\
        );

    \I__1759\ : InMux
    port map (
            O => \N__19124\,
            I => \N__19113\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19110\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__19116\,
            I => \N__19105\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__19113\,
            I => \N__19105\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__19110\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__19105\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__1753\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__19097\,
            I => \current_shift_inst.PI_CTRL.N_155\
        );

    \I__1751\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__1749\ : Span12Mux_h
    port map (
            O => \N__19088\,
            I => \N__19085\
        );

    \I__1748\ : Odrv12
    port map (
            O => \N__19085\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__1746\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__1744\ : Span4Mux_h
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__19070\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1742\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__19064\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__1740\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19058\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__19058\,
            I => \N__19055\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__19055\,
            I => \N__19052\
        );

    \I__1737\ : Span4Mux_v
    port map (
            O => \N__19052\,
            I => \N__19049\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__19049\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__1734\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__1732\ : Span4Mux_h
    port map (
            O => \N__19037\,
            I => \N__19034\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__19034\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__1729\ : InMux
    port map (
            O => \N__19028\,
            I => \N__19025\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__19025\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__1727\ : InMux
    port map (
            O => \N__19022\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1726\ : InMux
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__19016\,
            I => \N__19013\
        );

    \I__1724\ : Span4Mux_v
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__19010\,
            I => \N__19007\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__19007\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__1720\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__18992\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1716\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18986\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__18983\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__1713\ : InMux
    port map (
            O => \N__18980\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1712\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18974\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__18974\,
            I => \N__18971\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__18971\,
            I => \N__18968\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__18968\,
            I => \N__18965\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__18965\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__18962\,
            I => \N__18959\
        );

    \I__1706\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__18956\,
            I => \N__18953\
        );

    \I__1704\ : Span4Mux_h
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__18950\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__1701\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__18941\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__1699\ : InMux
    port map (
            O => \N__18938\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1698\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18932\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18929\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__18926\,
            I => \N__18923\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__18923\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__1692\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__18908\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1688\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__18899\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__1685\ : InMux
    port map (
            O => \N__18896\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1684\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__18881\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__1678\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__1675\ : Span4Mux_h
    port map (
            O => \N__18866\,
            I => \N__18863\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__18863\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__1672\ : InMux
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__18851\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__1669\ : InMux
    port map (
            O => \N__18848\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1668\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18840\
        );

    \I__1667\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18835\
        );

    \I__1666\ : InMux
    port map (
            O => \N__18843\,
            I => \N__18835\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__18840\,
            I => \N__18832\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__18835\,
            I => pwm_duty_input_4
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__18832\,
            I => pwm_duty_input_4
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__18827\,
            I => \N__18822\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__18826\,
            I => \N__18819\
        );

    \I__1660\ : InMux
    port map (
            O => \N__18825\,
            I => \N__18816\
        );

    \I__1659\ : InMux
    port map (
            O => \N__18822\,
            I => \N__18811\
        );

    \I__1658\ : InMux
    port map (
            O => \N__18819\,
            I => \N__18811\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__18816\,
            I => \N__18808\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__18811\,
            I => \N__18805\
        );

    \I__1655\ : Span4Mux_s1_h
    port map (
            O => \N__18808\,
            I => \N__18802\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__18805\,
            I => pwm_duty_input_3
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__18802\,
            I => pwm_duty_input_3
        );

    \I__1652\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18793\
        );

    \I__1651\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18790\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__18793\,
            I => \N__18787\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__18790\,
            I => pwm_duty_input_0
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__18787\,
            I => pwm_duty_input_0
        );

    \I__1647\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__18779\,
            I => \N__18775\
        );

    \I__1645\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18772\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__18775\,
            I => \N__18769\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__18772\,
            I => pwm_duty_input_1
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__18769\,
            I => pwm_duty_input_1
        );

    \I__1641\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__18761\,
            I => \N__18757\
        );

    \I__1639\ : InMux
    port map (
            O => \N__18760\,
            I => \N__18754\
        );

    \I__1638\ : Span4Mux_s1_h
    port map (
            O => \N__18757\,
            I => \N__18751\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__18754\,
            I => pwm_duty_input_2
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__18751\,
            I => pwm_duty_input_2
        );

    \I__1635\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__18743\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__18740\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__1631\ : InMux
    port map (
            O => \N__18734\,
            I => \N__18728\
        );

    \I__1630\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18728\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__18728\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__18725\,
            I => \current_shift_inst.PI_CTRL.N_31_cascade_\
        );

    \I__1627\ : InMux
    port map (
            O => \N__18722\,
            I => \N__18719\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__18716\,
            I => \current_shift_inst.PI_CTRL.N_149\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__18713\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\
        );

    \I__1623\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__18707\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__18704\,
            I => \current_shift_inst.PI_CTRL.N_27_cascade_\
        );

    \I__1620\ : InMux
    port map (
            O => \N__18701\,
            I => \N__18695\
        );

    \I__1619\ : InMux
    port map (
            O => \N__18700\,
            I => \N__18695\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__18692\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__18689\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\
        );

    \I__1615\ : InMux
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__18683\,
            I => \N_38_i_i\
        );

    \I__1613\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18677\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__18677\,
            I => \rgb_drv_RNOZ0\
        );

    \I__1611\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__18671\,
            I => \N__18668\
        );

    \I__1609\ : Span4Mux_h
    port map (
            O => \N__18668\,
            I => \N__18664\
        );

    \I__1608\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18661\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__18664\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__18661\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1605\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18653\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__18650\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \I__1602\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18638\
        );

    \I__1601\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18638\
        );

    \I__1600\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18638\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__18638\,
            I => \current_shift_inst.PI_CTRL.N_154\
        );

    \I__1598\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18632\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__18632\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__18629\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__18626\,
            I => \N__18622\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__18625\,
            I => \N__18619\
        );

    \I__1593\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18613\
        );

    \I__1592\ : InMux
    port map (
            O => \N__18619\,
            I => \N__18613\
        );

    \I__1591\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18610\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__18613\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__18610\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1588\ : InMux
    port map (
            O => \N__18605\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__1587\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18596\
        );

    \I__1586\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18596\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__18593\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__18590\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\
        );

    \I__1582\ : InMux
    port map (
            O => \N__18587\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__1581\ : InMux
    port map (
            O => \N__18584\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__1580\ : InMux
    port map (
            O => \N__18581\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__1579\ : InMux
    port map (
            O => \N__18578\,
            I => \bfn_1_15_0_\
        );

    \I__1578\ : IoInMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__1576\ : IoSpan4Mux
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__1575\ : Sp12to4
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__1574\ : Span12Mux_s6_v
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__1573\ : Span12Mux_h
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__1572\ : Odrv12
    port map (
            O => \N__18557\,
            I => \pll_inst.red_c_i\
        );

    \I__1571\ : InMux
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__1569\ : Odrv4
    port map (
            O => \N__18548\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1568\ : InMux
    port map (
            O => \N__18545\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1567\ : InMux
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__18536\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1564\ : InMux
    port map (
            O => \N__18533\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1563\ : InMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__18521\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1559\ : InMux
    port map (
            O => \N__18518\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1558\ : InMux
    port map (
            O => \N__18515\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__1557\ : IoInMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__1555\ : Span4Mux_s3_v
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__1554\ : Span4Mux_h
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__1553\ : Sp12to4
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__1552\ : Span12Mux_v
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__1551\ : Span12Mux_v
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__1550\ : Odrv12
    port map (
            O => \N__18491\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1549\ : IoInMux
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__1547\ : IoSpan4Mux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__1546\ : IoSpan4Mux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__1545\ : Odrv4
    port map (
            O => \N__18476\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_2_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_2_18_0_\
        );

    \IN_MUX_bfv_3_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_12_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_5_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_18_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_18_22_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_12_12_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18512\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18488\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__37628\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__23594\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_434_i_g\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__30617\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_432_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__39048\,
            CLKHFEN => \N__39068\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__39067\,
            RGB2PWM => \N__18686\,
            RGB1 => rgb_g_wire,
            CURREN => \N__38975\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__18680\,
            RGB0PWM => \N__47483\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__19541\,
            in1 => \N__18667\,
            in2 => \_gnd_net_\,
            in3 => \N__21358\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22253\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47876\,
            ce => 'H',
            sr => \N__47362\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__18618\,
            in1 => \N__21857\,
            in2 => \N__19130\,
            in3 => \N__18646\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47874\,
            ce => 'H',
            sr => \N__47386\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__18647\,
            in1 => \N__21845\,
            in2 => \N__18626\,
            in3 => \N__19129\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47874\,
            ce => 'H',
            sr => \N__47386\
        );

    \pwm_generator_inst.threshold_5_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20039\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47874\,
            ce => 'H',
            sr => \N__47386\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__18645\,
            in1 => \N__21866\,
            in2 => \N__18625\,
            in3 => \N__19128\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47874\,
            ce => 'H',
            sr => \N__47386\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101110"
        )
    port map (
            in0 => \N__21731\,
            in1 => \N__20257\,
            in2 => \N__20205\,
            in3 => \N__22243\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => 'H',
            sr => \N__47389\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101110"
        )
    port map (
            in0 => \N__21697\,
            in1 => \N__20258\,
            in2 => \N__20206\,
            in3 => \N__22244\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => 'H',
            sr => \N__47389\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111100001010"
        )
    port map (
            in0 => \N__20253\,
            in1 => \N__20191\,
            in2 => \N__22252\,
            in3 => \N__22030\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => 'H',
            sr => \N__47389\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__18710\,
            in1 => \N__21806\,
            in2 => \N__20204\,
            in3 => \N__18722\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => 'H',
            sr => \N__47389\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011111011"
        )
    port map (
            in0 => \N__21833\,
            in1 => \N__18635\,
            in2 => \N__20261\,
            in3 => \N__19123\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => 'H',
            sr => \N__47389\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101110"
        )
    port map (
            in0 => \N__21997\,
            in1 => \N__20259\,
            in2 => \N__20207\,
            in3 => \N__22248\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => 'H',
            sr => \N__47389\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__22242\,
            in1 => \N__20260\,
            in2 => \N__21761\,
            in3 => \N__20190\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47871\,
            ce => 'H',
            sr => \N__47395\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21246\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21220\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__47480\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19822\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18554\,
            in2 => \_gnd_net_\,
            in3 => \N__18545\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18542\,
            in2 => \_gnd_net_\,
            in3 => \N__18533\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18530\,
            in2 => \_gnd_net_\,
            in3 => \N__18518\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19067\,
            in2 => \_gnd_net_\,
            in3 => \N__18515\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38985\,
            in2 => \N__19031\,
            in3 => \N__18587\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18989\,
            in2 => \N__39055\,
            in3 => \N__18584\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38989\,
            in2 => \N__18947\,
            in3 => \N__18581\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18905\,
            in2 => \_gnd_net_\,
            in3 => \N__18578\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18860\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19367\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19325\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19283\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19244\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19220\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19196\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19172\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19145\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19568\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19466\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18605\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19424\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20093\,
            in2 => \_gnd_net_\,
            in3 => \N__18601\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__18602\,
            in1 => \N__21202\,
            in2 => \N__18590\,
            in3 => \N__20081\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18700\,
            in2 => \_gnd_net_\,
            in3 => \N__20072\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__18701\,
            in1 => \N__21203\,
            in2 => \N__18689\,
            in3 => \N__20060\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20476\,
            in2 => \_gnd_net_\,
            in3 => \N__20449\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_0_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__47481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34159\,
            lcout => \N_38_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__47482\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34163\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__18674\,
            in1 => \N__19540\,
            in2 => \N__21379\,
            in3 => \N__18656\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__22240\,
            in1 => \_gnd_net_\,
            in2 => \N__18737\,
            in3 => \N__20233\,
            lcout => \current_shift_inst.PI_CTRL.N_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__21797\,
            in1 => \N__22239\,
            in2 => \_gnd_net_\,
            in3 => \N__18733\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010000"
        )
    port map (
            in0 => \N__21831\,
            in1 => \N__20234\,
            in2 => \N__18629\,
            in3 => \N__19124\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101011"
        )
    port map (
            in0 => \N__19928\,
            in1 => \N__18844\,
            in2 => \N__18826\,
            in3 => \N__18746\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__20045\,
            in1 => \N__18843\,
            in2 => \N__18827\,
            in3 => \N__20290\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__18796\,
            in1 => \N__18778\,
            in2 => \_gnd_net_\,
            in3 => \N__18760\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__21996\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21756\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22029\,
            in1 => \N__21696\,
            in2 => \N__18740\,
            in3 => \N__21730\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => \current_shift_inst.PI_CTRL.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__21805\,
            in1 => \N__22241\,
            in2 => \N__18725\,
            in3 => \N__20235\,
            lcout => \current_shift_inst.PI_CTRL.N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22001\,
            in2 => \_gnd_net_\,
            in3 => \N__21729\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22031\,
            in1 => \N__21698\,
            in2 => \N__18713\,
            in3 => \N__21757\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => \current_shift_inst.PI_CTRL.N_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__22215\,
            in1 => \N__19100\,
            in2 => \N__18704\,
            in3 => \N__20172\,
            lcout => \current_shift_inst.PI_CTRL.N_153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21801\,
            in2 => \_gnd_net_\,
            in3 => \N__21832\,
            lcout => \current_shift_inst.PI_CTRL.N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19094\,
            in2 => \N__19082\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19061\,
            in2 => \N__19046\,
            in3 => \N__19022\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19019\,
            in2 => \N__19004\,
            in3 => \N__18980\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18977\,
            in2 => \N__18962\,
            in3 => \N__18938\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18935\,
            in2 => \N__18920\,
            in3 => \N__18896\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18893\,
            in2 => \N__18878\,
            in3 => \N__18848\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19394\,
            in2 => \N__19382\,
            in3 => \N__19358\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19355\,
            in2 => \N__19340\,
            in3 => \N__19313\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19310\,
            in2 => \N__19298\,
            in3 => \N__19277\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19274\,
            in2 => \N__19259\,
            in3 => \N__19238\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19235\,
            in2 => \N__19535\,
            in3 => \N__19214\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19211\,
            in2 => \N__19537\,
            in3 => \N__19190\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19187\,
            in2 => \N__19536\,
            in3 => \N__19163\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19160\,
            in2 => \N__19538\,
            in3 => \N__19133\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19525\,
            in2 => \N__19583\,
            in3 => \N__19559\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19556\,
            in2 => \N__19539\,
            in3 => \N__19454\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19451\,
            in1 => \N__19439\,
            in2 => \_gnd_net_\,
            in3 => \N__19427\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__19784\,
            in1 => \N__19423\,
            in2 => \N__19409\,
            in3 => \N__19801\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20658\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19405\,
            in2 => \_gnd_net_\,
            in3 => \N__20119\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__19406\,
            in1 => \N__21169\,
            in2 => \N__19397\,
            in3 => \N__20105\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19738\,
            in2 => \_gnd_net_\,
            in3 => \N__19768\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19739\,
            in1 => \N__19754\,
            in2 => \N__19730\,
            in3 => \N__21168\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19712\,
            in2 => \_gnd_net_\,
            in3 => \N__19727\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19691\,
            in2 => \_gnd_net_\,
            in3 => \N__19706\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19670\,
            in2 => \_gnd_net_\,
            in3 => \N__19685\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19649\,
            in2 => \_gnd_net_\,
            in3 => \N__19664\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19628\,
            in2 => \_gnd_net_\,
            in3 => \N__19643\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19607\,
            in2 => \_gnd_net_\,
            in3 => \N__19622\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19589\,
            in2 => \_gnd_net_\,
            in3 => \N__19601\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19880\,
            in2 => \_gnd_net_\,
            in3 => \N__19895\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19859\,
            in2 => \_gnd_net_\,
            in3 => \N__19874\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19838\,
            in2 => \_gnd_net_\,
            in3 => \N__19853\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20445\,
            in2 => \_gnd_net_\,
            in3 => \N__19832\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__21176\,
            in1 => \N__19829\,
            in2 => \_gnd_net_\,
            in3 => \N__19805\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19800\,
            in2 => \_gnd_net_\,
            in3 => \N__19775\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21253\,
            in2 => \_gnd_net_\,
            in3 => \N__19772\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19769\,
            in2 => \_gnd_net_\,
            in3 => \N__19742\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20120\,
            in2 => \_gnd_net_\,
            in3 => \N__20096\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20092\,
            in2 => \_gnd_net_\,
            in3 => \N__20075\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_18_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20071\,
            in2 => \_gnd_net_\,
            in3 => \N__20054\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20662\,
            in2 => \_gnd_net_\,
            in3 => \N__20051\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20048\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19922\,
            in1 => \N__19999\,
            in2 => \N__19963\,
            in3 => \N__20030\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__21486\,
            in1 => \N__20756\,
            in2 => \N__21439\,
            in3 => \N__21554\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47872\,
            ce => 'H',
            sr => \N__47371\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__20026\,
            in1 => \N__20000\,
            in2 => \N__19964\,
            in3 => \N__20270\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__19921\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20294\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20213\,
            in1 => \N__21959\,
            in2 => \N__21941\,
            in3 => \N__20807\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20903\,
            in1 => \N__20801\,
            in2 => \N__20264\,
            in3 => \N__20600\,
            lcout => \current_shift_inst.PI_CTRL.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22142\,
            in2 => \_gnd_net_\,
            in3 => \N__22160\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20771\,
            in1 => \N__20813\,
            in2 => \N__20795\,
            in3 => \N__20783\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20312\,
            in2 => \N__20156\,
            in3 => \N__20878\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_3_12_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20856\,
            in1 => \N__20303\,
            in2 => \N__20147\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20135\,
            in2 => \N__20915\,
            in3 => \N__20836\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21656\,
            in2 => \N__20129\,
            in3 => \N__21111\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20399\,
            in2 => \N__20498\,
            in3 => \N__21090\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20378\,
            in2 => \N__20393\,
            in3 => \N__21069\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20486\,
            in2 => \N__20372\,
            in3 => \N__21048\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21027\,
            in1 => \N__20588\,
            in2 => \N__20363\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21614\,
            in2 => \N__20354\,
            in3 => \N__21006\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21665\,
            in2 => \N__20345\,
            in3 => \N__20934\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20336\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47860\,
            ce => 'H',
            sr => \N__47396\
        );

    \pwm_generator_inst.threshold_0_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20417\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => 'H',
            sr => \N__47401\
        );

    \pwm_generator_inst.threshold_1_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20570\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => 'H',
            sr => \N__47401\
        );

    \pwm_generator_inst.threshold_4_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20579\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => 'H',
            sr => \N__47401\
        );

    \pwm_generator_inst.threshold_6_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20408\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => 'H',
            sr => \N__47401\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20477\,
            in1 => \N__20453\,
            in2 => \N__20429\,
            in3 => \N__21167\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__27162\,
            in1 => \N__27347\,
            in2 => \N__27431\,
            in3 => \N__24461\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__24365\,
            sr => \N__47407\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27344\,
            in1 => \N__27163\,
            in2 => \N__27539\,
            in3 => \N__24469\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__24365\,
            sr => \N__47407\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27161\,
            in1 => \N__27346\,
            in2 => \N__31256\,
            in3 => \N__24460\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__24365\,
            sr => \N__47407\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27345\,
            in1 => \N__27164\,
            in2 => \N__27470\,
            in3 => \N__24470\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__24365\,
            sr => \N__47407\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__21582\,
            in1 => \N__20552\,
            in2 => \N__21434\,
            in3 => \N__21512\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__47414\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__21515\,
            in1 => \N__20732\,
            in2 => \N__21437\,
            in3 => \N__21585\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__47414\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__21516\,
            in1 => \N__20714\,
            in2 => \N__21438\,
            in3 => \N__21586\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__47414\
        );

    \pwm_generator_inst.threshold_7_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20594\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__47414\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__21584\,
            in1 => \N__20507\,
            in2 => \N__21435\,
            in3 => \N__21514\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__47414\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__21513\,
            in1 => \N__20540\,
            in2 => \N__21436\,
            in3 => \N__21583\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__47414\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20561\,
            in2 => \N__21208\,
            in3 => \N__21201\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20546\,
            in2 => \_gnd_net_\,
            in3 => \N__20534\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20531\,
            in2 => \_gnd_net_\,
            in3 => \N__20522\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21119\,
            in2 => \_gnd_net_\,
            in3 => \N__20519\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20516\,
            in2 => \_gnd_net_\,
            in3 => \N__20501\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20765\,
            in2 => \_gnd_net_\,
            in3 => \N__20744\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20741\,
            in2 => \_gnd_net_\,
            in3 => \N__20726\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20723\,
            in2 => \_gnd_net_\,
            in3 => \N__20708\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20633\,
            in2 => \_gnd_net_\,
            in3 => \N__20705\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__20702\,
            in1 => \N__20690\,
            in2 => \N__21209\,
            in3 => \N__20684\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__20681\,
            in1 => \N__21204\,
            in2 => \N__20663\,
            in3 => \N__20639\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20627\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22280\,
            in1 => \N__22334\,
            in2 => \N__22316\,
            in3 => \N__20777\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21934\,
            in2 => \_gnd_net_\,
            in3 => \N__21970\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21955\,
            in1 => \N__22312\,
            in2 => \N__20816\,
            in3 => \N__20897\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22298\,
            in1 => \N__21971\,
            in2 => \N__22178\,
            in3 => \N__21890\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21920\,
            in1 => \N__22067\,
            in2 => \N__22052\,
            in3 => \N__21905\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22330\,
            in1 => \N__22138\,
            in2 => \N__22276\,
            in3 => \N__22156\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22174\,
            in2 => \_gnd_net_\,
            in3 => \N__21889\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22079\,
            in1 => \N__22345\,
            in2 => \N__20786\,
            in3 => \N__22360\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22096\,
            in2 => \_gnd_net_\,
            in3 => \N__22078\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22123\,
            in1 => \N__21904\,
            in2 => \N__22112\,
            in3 => \N__21919\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22361\,
            in1 => \N__22111\,
            in2 => \N__22349\,
            in3 => \N__22124\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22294\,
            in1 => \N__22066\,
            in2 => \N__22097\,
            in3 => \N__22045\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__20835\,
            in1 => \N__20877\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__21091\,
            in1 => \N__20857\,
            in2 => \N__20891\,
            in3 => \N__21112\,
            lcout => \pwm_generator_inst.un1_counterlt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20936\,
            in1 => \N__21008\,
            in2 => \_gnd_net_\,
            in3 => \N__21028\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21050\,
            in1 => \N__21071\,
            in2 => \N__20888\,
            in3 => \N__20885\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20981\,
            in1 => \N__20879\,
            in2 => \_gnd_net_\,
            in3 => \N__20861\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__47390\
        );

    \pwm_generator_inst.counter_1_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20966\,
            in1 => \N__20858\,
            in2 => \_gnd_net_\,
            in3 => \N__20840\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__47390\
        );

    \pwm_generator_inst.counter_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20982\,
            in1 => \N__20837\,
            in2 => \_gnd_net_\,
            in3 => \N__20819\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__47390\
        );

    \pwm_generator_inst.counter_3_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20967\,
            in1 => \N__21113\,
            in2 => \_gnd_net_\,
            in3 => \N__21095\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__47390\
        );

    \pwm_generator_inst.counter_4_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20983\,
            in1 => \N__21092\,
            in2 => \_gnd_net_\,
            in3 => \N__21074\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__47390\
        );

    \pwm_generator_inst.counter_5_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20968\,
            in1 => \N__21070\,
            in2 => \_gnd_net_\,
            in3 => \N__21053\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__47390\
        );

    \pwm_generator_inst.counter_6_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20984\,
            in1 => \N__21049\,
            in2 => \_gnd_net_\,
            in3 => \N__21032\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__47390\
        );

    \pwm_generator_inst.counter_7_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20969\,
            in1 => \N__21029\,
            in2 => \_gnd_net_\,
            in3 => \N__21011\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__47390\
        );

    \pwm_generator_inst.counter_8_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20980\,
            in1 => \N__21007\,
            in2 => \_gnd_net_\,
            in3 => \N__20987\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__47840\,
            ce => 'H',
            sr => \N__47397\
        );

    \pwm_generator_inst.counter_9_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__20935\,
            in1 => \N__20979\,
            in2 => \_gnd_net_\,
            in3 => \N__20939\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47840\,
            ce => 'H',
            sr => \N__47397\
        );

    \pwm_generator_inst.threshold_2_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21635\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47840\,
            ce => 'H',
            sr => \N__47397\
        );

    \pwm_generator_inst.threshold_9_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21275\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47832\,
            ce => 'H',
            sr => \N__47402\
        );

    \pwm_generator_inst.threshold_3_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21620\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47826\,
            ce => 'H',
            sr => \N__47408\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__21589\,
            in1 => \N__21464\,
            in2 => \N__21644\,
            in3 => \N__21527\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47826\,
            ce => 'H',
            sr => \N__47408\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__21528\,
            in1 => \N__21590\,
            in2 => \N__21470\,
            in3 => \N__21626\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47826\,
            ce => 'H',
            sr => \N__47408\
        );

    \pwm_generator_inst.threshold_8_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21596\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47826\,
            ce => 'H',
            sr => \N__47408\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__21587\,
            in1 => \N__21602\,
            in2 => \N__21469\,
            in3 => \N__21529\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => 'H',
            sr => \N__47415\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__21588\,
            in1 => \N__21530\,
            in2 => \N__21468\,
            in3 => \N__21281\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => 'H',
            sr => \N__47415\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__21266\,
            in1 => \N__21257\,
            in2 => \N__21230\,
            in3 => \N__21197\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21875\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28358\,
            in2 => \N__23579\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28337\,
            in2 => \N__30569\,
            in3 => \N__21848\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26176\,
            in2 => \N__30803\,
            in3 => \N__21836\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22478\,
            in2 => \N__25714\,
            in3 => \N__21809\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25754\,
            in2 => \N__28604\,
            in3 => \N__21764\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25795\,
            in2 => \N__28589\,
            in3 => \N__21734\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28426\,
            in2 => \N__22406\,
            in3 => \N__21701\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28346\,
            in2 => \N__22769\,
            in3 => \N__21668\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22499\,
            in2 => \N__30782\,
            in3 => \N__22004\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__47865\,
            ce => 'H',
            sr => \N__47363\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25948\,
            in2 => \N__22490\,
            in3 => \N__21974\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__47865\,
            ce => 'H',
            sr => \N__47363\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22967\,
            in2 => \N__26015\,
            in3 => \N__21962\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__47865\,
            ce => 'H',
            sr => \N__47363\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22466\,
            in2 => \N__25510\,
            in3 => \N__21944\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__47865\,
            ce => 'H',
            sr => \N__47363\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22925\,
            in2 => \N__28490\,
            in3 => \N__21923\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__47865\,
            ce => 'H',
            sr => \N__47363\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40546\,
            in2 => \N__22951\,
            in3 => \N__21908\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__47865\,
            ce => 'H',
            sr => \N__47363\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22929\,
            in2 => \N__25565\,
            in3 => \N__21893\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__47865\,
            ce => 'H',
            sr => \N__47363\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24047\,
            in2 => \N__22952\,
            in3 => \N__21878\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__47865\,
            ce => 'H',
            sr => \N__47363\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22892\,
            in2 => \N__25381\,
            in3 => \N__22163\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47372\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25855\,
            in2 => \N__22933\,
            in3 => \N__22145\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47372\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22896\,
            in2 => \N__25907\,
            in3 => \N__22127\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47372\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27599\,
            in2 => \N__22934\,
            in3 => \N__22115\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47372\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22900\,
            in2 => \N__26237\,
            in3 => \N__22100\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47372\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30697\,
            in2 => \N__22935\,
            in3 => \N__22082\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47372\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22904\,
            in2 => \N__26072\,
            in3 => \N__22070\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47372\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26359\,
            in2 => \N__22936\,
            in3 => \N__22055\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47372\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22937\,
            in2 => \N__30500\,
            in3 => \N__22034\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__47849\,
            ce => 'H',
            sr => \N__47378\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26300\,
            in2 => \N__22953\,
            in3 => \N__22352\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__47849\,
            ce => 'H',
            sr => \N__47378\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22941\,
            in2 => \N__26126\,
            in3 => \N__22337\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__47849\,
            ce => 'H',
            sr => \N__47378\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29272\,
            in2 => \N__22954\,
            in3 => \N__22319\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__47849\,
            ce => 'H',
            sr => \N__47378\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22945\,
            in2 => \N__24098\,
            in3 => \N__22301\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__47849\,
            ce => 'H',
            sr => \N__47378\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24135\,
            in2 => \N__22955\,
            in3 => \N__22283\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__47849\,
            ce => 'H',
            sr => \N__47378\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22949\,
            in2 => \N__40613\,
            in3 => \N__22259\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__47849\,
            ce => 'H',
            sr => \N__47378\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22950\,
            in1 => \N__28305\,
            in2 => \_gnd_net_\,
            in3 => \N__22256\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47849\,
            ce => 'H',
            sr => \N__47378\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22190\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26364\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25890\,
            in1 => \N__25840\,
            in2 => \N__24041\,
            in3 => \N__26226\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26363\,
            in1 => \N__25380\,
            in2 => \N__26014\,
            in3 => \N__24136\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25379\,
            in1 => \N__26006\,
            in2 => \N__24140\,
            in3 => \N__26365\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22433\,
            in1 => \N__22814\,
            in2 => \N__25406\,
            in3 => \N__22391\,
            lcout => \current_shift_inst.PI_CTRL.N_74_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__26054\,
            in1 => \N__25509\,
            in2 => \_gnd_net_\,
            in3 => \N__22382\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25421\,
            in1 => \N__22376\,
            in2 => \N__22370\,
            in3 => \N__22412\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__22427\,
            in1 => \N__25750\,
            in2 => \N__22367\,
            in3 => \N__22451\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__25655\,
            in1 => \N__22439\,
            in2 => \N__22364\,
            in3 => \N__22831\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26005\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__22846\,
            in1 => \_gnd_net_\,
            in2 => \N__25511\,
            in3 => \N__28317\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30475\,
            in1 => \N__30679\,
            in2 => \N__27596\,
            in3 => \N__26102\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26101\,
            in1 => \N__24096\,
            in2 => \N__29271\,
            in3 => \N__26279\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__25713\,
            in1 => \N__30568\,
            in2 => \N__26180\,
            in3 => \N__23571\,
            lcout => \current_shift_inst.PI_CTRL.N_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25889\,
            in1 => \N__25842\,
            in2 => \N__24040\,
            in3 => \N__26215\,
            lcout => \current_shift_inst.PI_CTRL.N_74_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29263\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24097\,
            in2 => \_gnd_net_\,
            in3 => \N__26278\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40601\,
            in1 => \N__29264\,
            in2 => \N__22421\,
            in3 => \N__22418\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30869\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47850\,
            ce => 'H',
            sr => \N__47341\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31094\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47850\,
            ce => 'H',
            sr => \N__47341\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31061\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47850\,
            ce => 'H',
            sr => \N__47341\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30947\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47850\,
            ce => 'H',
            sr => \N__47341\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31133\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47850\,
            ce => 'H',
            sr => \N__47341\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22761\,
            in2 => \_gnd_net_\,
            in3 => \N__25785\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22762\,
            in1 => \N__30768\,
            in2 => \N__28419\,
            in3 => \N__25935\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25934\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__28269\,
            in1 => \N__23882\,
            in2 => \N__28152\,
            in3 => \N__27977\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47841\,
            ce => 'H',
            sr => \N__47353\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__25936\,
            in1 => \N__22457\,
            in2 => \N__30781\,
            in3 => \N__28415\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23572\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33678\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28839\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__28974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33677\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23343\,
            in1 => \N__23441\,
            in2 => \N__22553\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23092\,
            in1 => \N__23387\,
            in2 => \N__22544\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23453\,
            in2 => \N__22535\,
            in3 => \N__23074\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23375\,
            in2 => \N__22526\,
            in3 => \N__23059\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23044\,
            in1 => \N__23477\,
            in2 => \N__22517\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23399\,
            in2 => \N__22508\,
            in3 => \N__23029\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24377\,
            in2 => \N__22670\,
            in3 => \N__23014\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23465\,
            in2 => \N__22661\,
            in3 => \N__22999\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22981\,
            in1 => \N__24245\,
            in2 => \N__22652\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22643\,
            in2 => \N__22631\,
            in3 => \N__23227\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22622\,
            in2 => \N__22610\,
            in3 => \N__23212\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22601\,
            in2 => \N__22589\,
            in3 => \N__23197\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23182\,
            in1 => \N__22580\,
            in2 => \N__24236\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22574\,
            in2 => \N__22562\,
            in3 => \N__23167\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24179\,
            in2 => \N__22721\,
            in3 => \N__23152\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23137\,
            in1 => \N__24188\,
            in2 => \N__22709\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23122\,
            in1 => \N__24200\,
            in2 => \N__22700\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24212\,
            in2 => \N__22691\,
            in3 => \N__23107\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24224\,
            in2 => \N__22682\,
            in3 => \N__23359\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22673\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_0_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36284\,
            in1 => \N__36252\,
            in2 => \_gnd_net_\,
            in3 => \N__23300\,
            lcout => \phase_controller_inst1.stoper_hc.running_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000101110"
        )
    port map (
            in0 => \N__23264\,
            in1 => \N__23249\,
            in2 => \N__36300\,
            in3 => \N__23321\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47809\,
            ce => 'H',
            sr => \N__47391\
        );

    \phase_controller_inst2.start_timer_hc_RNO_1_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32419\,
            in2 => \_gnd_net_\,
            in3 => \N__32067\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__34827\,
            in1 => \N__22730\,
            in2 => \N__22733\,
            in3 => \N__27738\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47809\,
            ce => 'H',
            sr => \N__47391\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32138\,
            in2 => \_gnd_net_\,
            in3 => \N__32112\,
            lcout => \phase_controller_inst2.start_timer_hc_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_2_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__32139\,
            in1 => \N__32113\,
            in2 => \N__32074\,
            in3 => \N__32420\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47809\,
            ce => 'H',
            sr => \N__47391\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36253\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47809\,
            ce => 'H',
            sr => \N__47391\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__22793\,
            in1 => \N__27015\,
            in2 => \N__22808\,
            in3 => \N__24801\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => 'H',
            sr => \N__47403\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22792\,
            in2 => \_gnd_net_\,
            in3 => \N__22804\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__34598\,
            in1 => \N__34625\,
            in2 => \N__35742\,
            in3 => \N__42102\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => 'H',
            sr => \N__47403\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__27698\,
            in1 => \N__32111\,
            in2 => \N__27750\,
            in3 => \N__27653\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__47409\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__27666\,
            in1 => \N__27696\,
            in2 => \_gnd_net_\,
            in3 => \N__27739\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.running_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001011100"
        )
    port map (
            in0 => \N__27699\,
            in1 => \N__27667\,
            in2 => \N__22724\,
            in3 => \N__27761\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__47409\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27743\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__47409\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27697\,
            in2 => \_gnd_net_\,
            in3 => \N__27782\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22796\,
            in3 => \N__22791\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27705\,
            in2 => \_gnd_net_\,
            in3 => \N__27749\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22778\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25841\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__22752\,
            in1 => \N__33774\,
            in2 => \N__31132\,
            in3 => \N__28712\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22751\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__28316\,
            in1 => \N__28143\,
            in2 => \N__27979\,
            in3 => \N__23675\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47862\,
            ce => 'H',
            sr => \N__47330\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110100001100"
        )
    port map (
            in0 => \N__23846\,
            in1 => \N__28314\,
            in2 => \N__28165\,
            in3 => \N__27935\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47862\,
            ce => 'H',
            sr => \N__47330\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__28145\,
            in1 => \N__23807\,
            in2 => \N__27980\,
            in3 => \N__28315\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47862\,
            ce => 'H',
            sr => \N__47330\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__28313\,
            in1 => \N__28144\,
            in2 => \N__27978\,
            in3 => \N__23786\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47862\,
            ce => 'H',
            sr => \N__47330\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__25775\,
            in1 => \N__31057\,
            in2 => \N__33776\,
            in3 => \N__28742\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25774\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__28002\,
            in1 => \N__28304\,
            in2 => \N__23726\,
            in3 => \N__28100\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47851\,
            ce => 'H',
            sr => \N__47333\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28300\,
            in1 => \N__28003\,
            in2 => \N__28148\,
            in3 => \N__23774\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47851\,
            ce => 'H',
            sr => \N__47333\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28000\,
            in1 => \N__28302\,
            in2 => \N__23756\,
            in3 => \N__28098\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47851\,
            ce => 'H',
            sr => \N__47333\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28301\,
            in1 => \N__28004\,
            in2 => \N__28149\,
            in3 => \N__23981\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47851\,
            ce => 'H',
            sr => \N__47333\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28001\,
            in1 => \N__28303\,
            in2 => \N__23969\,
            in3 => \N__28099\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47851\,
            ce => 'H',
            sr => \N__47333\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30476\,
            in1 => \N__30680\,
            in2 => \N__27597\,
            in3 => \N__26053\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22847\,
            in1 => \N__25490\,
            in2 => \N__22835\,
            in3 => \N__25654\,
            lcout => \current_shift_inst.PI_CTRL.N_103\,
            ltout => \current_shift_inst.PI_CTRL.N_103_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28296\,
            in1 => \N__27952\,
            in2 => \N__22817\,
            in3 => \N__23606\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47842\,
            ce => 'H',
            sr => \N__47335\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25489\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28297\,
            in1 => \N__27953\,
            in2 => \N__28160\,
            in3 => \N__23936\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47842\,
            ce => 'H',
            sr => \N__47335\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__27951\,
            in1 => \N__28299\,
            in2 => \N__23927\,
            in3 => \N__28129\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47842\,
            ce => 'H',
            sr => \N__47335\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28298\,
            in1 => \N__27954\,
            in2 => \N__28161\,
            in3 => \N__23903\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47842\,
            ce => 'H',
            sr => \N__47335\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28265\,
            in1 => \N__27956\,
            in2 => \N__28147\,
            in3 => \N__23945\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => 'H',
            sr => \N__47342\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__27955\,
            in1 => \N__28266\,
            in2 => \N__28150\,
            in3 => \N__24158\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => 'H',
            sr => \N__47342\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__28264\,
            in1 => \N__23825\,
            in2 => \N__28146\,
            in3 => \N__27960\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => 'H',
            sr => \N__47342\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31028\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => 'H',
            sr => \N__47342\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33773\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => 'H',
            sr => \N__47342\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__23702\,
            in1 => \N__28267\,
            in2 => \N__28151\,
            in3 => \N__27961\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => 'H',
            sr => \N__47342\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__28101\,
            in1 => \N__28268\,
            in2 => \N__27996\,
            in3 => \N__23648\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => 'H',
            sr => \N__47342\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28408\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28261\,
            in1 => \N__27983\,
            in2 => \N__28163\,
            in3 => \N__23870\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47827\,
            ce => 'H',
            sr => \N__47354\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__27981\,
            in1 => \N__28263\,
            in2 => \N__24170\,
            in3 => \N__28139\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47827\,
            ce => 'H',
            sr => \N__47354\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28262\,
            in1 => \N__27984\,
            in2 => \N__28164\,
            in3 => \N__24146\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47827\,
            ce => 'H',
            sr => \N__47354\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__28260\,
            in1 => \N__27982\,
            in2 => \N__28162\,
            in3 => \N__23624\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47827\,
            ce => 'H',
            sr => \N__47354\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23309\,
            in2 => \N__23348\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24352\,
            in1 => \N__23093\,
            in2 => \_gnd_net_\,
            in3 => \N__23081\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__47821\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__24323\,
            in1 => \N__23273\,
            in2 => \N__23078\,
            in3 => \N__23063\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__47821\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24353\,
            in1 => \N__23060\,
            in2 => \_gnd_net_\,
            in3 => \N__23048\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__47821\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24324\,
            in1 => \N__23045\,
            in2 => \_gnd_net_\,
            in3 => \N__23033\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__47821\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24354\,
            in1 => \N__23030\,
            in2 => \_gnd_net_\,
            in3 => \N__23018\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__47821\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24325\,
            in1 => \N__23015\,
            in2 => \_gnd_net_\,
            in3 => \N__23003\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__47821\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24355\,
            in1 => \N__23000\,
            in2 => \_gnd_net_\,
            in3 => \N__22985\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__47821\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24364\,
            in1 => \N__22982\,
            in2 => \_gnd_net_\,
            in3 => \N__22970\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__47816\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24326\,
            in1 => \N__23228\,
            in2 => \_gnd_net_\,
            in3 => \N__23216\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__47816\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24361\,
            in1 => \N__23213\,
            in2 => \_gnd_net_\,
            in3 => \N__23201\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__47816\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24327\,
            in1 => \N__23198\,
            in2 => \_gnd_net_\,
            in3 => \N__23186\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__47816\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24362\,
            in1 => \N__23183\,
            in2 => \_gnd_net_\,
            in3 => \N__23171\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__47816\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24328\,
            in1 => \N__23168\,
            in2 => \_gnd_net_\,
            in3 => \N__23156\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__47816\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24363\,
            in1 => \N__23153\,
            in2 => \_gnd_net_\,
            in3 => \N__23141\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__47816\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24329\,
            in1 => \N__23138\,
            in2 => \_gnd_net_\,
            in3 => \N__23126\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__47816\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24330\,
            in1 => \N__23123\,
            in2 => \_gnd_net_\,
            in3 => \N__23111\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__47810\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24360\,
            in1 => \N__23108\,
            in2 => \_gnd_net_\,
            in3 => \N__23096\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__47810\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24331\,
            in1 => \N__23360\,
            in2 => \_gnd_net_\,
            in3 => \N__23363\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47810\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__23248\,
            in1 => \N__23288\,
            in2 => \N__23347\,
            in3 => \N__24332\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47810\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__24870\,
            in1 => \N__26550\,
            in2 => \N__24953\,
            in3 => \N__24406\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47803\,
            ce => \N__27021\,
            sr => \N__47387\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__23263\,
            in1 => \N__36241\,
            in2 => \N__36293\,
            in3 => \N__23320\,
            lcout => \phase_controller_inst1.stoper_hc.un1_start_latched2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23246\,
            in2 => \_gnd_net_\,
            in3 => \N__23287\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNI5B6O_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__36240\,
            in1 => \N__36280\,
            in2 => \_gnd_net_\,
            in3 => \N__23299\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTI1_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23276\,
            in3 => \N__23247\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNIQVTIZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__36239\,
            in1 => \N__23262\,
            in2 => \_gnd_net_\,
            in3 => \N__36279\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__24941\,
            in1 => \N__24871\,
            in2 => \N__24581\,
            in3 => \N__27297\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47799\,
            ce => \N__27020\,
            sr => \N__47392\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27293\,
            in1 => \N__26860\,
            in2 => \_gnd_net_\,
            in3 => \N__24943\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47799\,
            ce => \N__27020\,
            sr => \N__47392\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27294\,
            in1 => \N__26831\,
            in2 => \_gnd_net_\,
            in3 => \N__24944\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47799\,
            ce => \N__27020\,
            sr => \N__47392\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__27149\,
            in1 => \N__27292\,
            in2 => \_gnd_net_\,
            in3 => \N__33940\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47799\,
            ce => \N__27020\,
            sr => \N__47392\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__27295\,
            in1 => \N__24863\,
            in2 => \N__26798\,
            in3 => \N__24942\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47799\,
            ce => \N__27020\,
            sr => \N__47392\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__26646\,
            in1 => \N__27150\,
            in2 => \_gnd_net_\,
            in3 => \N__27296\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47799\,
            ce => \N__27020\,
            sr => \N__47392\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__24518\,
            in1 => \N__24535\,
            in2 => \N__24875\,
            in3 => \N__24388\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47799\,
            ce => \N__27020\,
            sr => \N__47392\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__24580\,
            in1 => \N__24869\,
            in2 => \N__24951\,
            in3 => \N__27350\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47794\,
            ce => \N__24356\,
            sr => \N__47398\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__24867\,
            in1 => \N__24497\,
            in2 => \N__27359\,
            in3 => \N__24938\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47794\,
            ce => \N__24356\,
            sr => \N__47398\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__24866\,
            in1 => \N__26702\,
            in2 => \N__24950\,
            in3 => \N__27349\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47794\,
            ce => \N__24356\,
            sr => \N__47398\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__27354\,
            in1 => \N__24940\,
            in2 => \N__26797\,
            in3 => \N__24865\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47794\,
            ce => \N__24356\,
            sr => \N__47398\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27348\,
            in2 => \N__24952\,
            in3 => \N__26827\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47794\,
            ce => \N__24356\,
            sr => \N__47398\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__24868\,
            in1 => \N__24939\,
            in2 => \N__24407\,
            in3 => \N__26554\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47794\,
            ce => \N__24356\,
            sr => \N__47398\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__24864\,
            in1 => \N__24389\,
            in2 => \N__24536\,
            in3 => \N__24517\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47794\,
            ce => \N__24356\,
            sr => \N__47398\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__40484\,
            in1 => \N__44077\,
            in2 => \_gnd_net_\,
            in3 => \N__40835\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23429\,
            in2 => \N__24805\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26960\,
            in1 => \N__24764\,
            in2 => \_gnd_net_\,
            in3 => \N__23423\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__47788\,
            ce => 'H',
            sr => \N__47404\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__26964\,
            in1 => \N__24743\,
            in2 => \N__23420\,
            in3 => \N__23408\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__47788\,
            ce => 'H',
            sr => \N__47404\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26961\,
            in1 => \N__24706\,
            in2 => \_gnd_net_\,
            in3 => \N__23405\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__47788\,
            ce => 'H',
            sr => \N__47404\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26965\,
            in1 => \N__24665\,
            in2 => \_gnd_net_\,
            in3 => \N__23402\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__47788\,
            ce => 'H',
            sr => \N__47404\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26962\,
            in1 => \N__24644\,
            in2 => \_gnd_net_\,
            in3 => \N__23504\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__47788\,
            ce => 'H',
            sr => \N__47404\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26966\,
            in1 => \N__24602\,
            in2 => \_gnd_net_\,
            in3 => \N__23501\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__47788\,
            ce => 'H',
            sr => \N__47404\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26963\,
            in1 => \N__25159\,
            in2 => \_gnd_net_\,
            in3 => \N__23498\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__47788\,
            ce => 'H',
            sr => \N__47404\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27009\,
            in1 => \N__25127\,
            in2 => \_gnd_net_\,
            in3 => \N__23495\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__47784\,
            ce => 'H',
            sr => \N__47410\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26953\,
            in1 => \N__25100\,
            in2 => \_gnd_net_\,
            in3 => \N__23492\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__47784\,
            ce => 'H',
            sr => \N__47410\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27006\,
            in1 => \N__25067\,
            in2 => \_gnd_net_\,
            in3 => \N__23489\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__47784\,
            ce => 'H',
            sr => \N__47410\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26954\,
            in1 => \N__25034\,
            in2 => \_gnd_net_\,
            in3 => \N__23486\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__47784\,
            ce => 'H',
            sr => \N__47410\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27007\,
            in1 => \N__25007\,
            in2 => \_gnd_net_\,
            in3 => \N__23483\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__47784\,
            ce => 'H',
            sr => \N__47410\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26955\,
            in1 => \N__24974\,
            in2 => \_gnd_net_\,
            in3 => \N__23480\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__47784\,
            ce => 'H',
            sr => \N__47410\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27008\,
            in1 => \N__25325\,
            in2 => \_gnd_net_\,
            in3 => \N__23519\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__47784\,
            ce => 'H',
            sr => \N__47410\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26956\,
            in1 => \N__25298\,
            in2 => \_gnd_net_\,
            in3 => \N__23516\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__47784\,
            ce => 'H',
            sr => \N__47410\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26957\,
            in1 => \N__25277\,
            in2 => \_gnd_net_\,
            in3 => \N__23513\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__47779\,
            ce => 'H',
            sr => \N__47416\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26959\,
            in1 => \N__25244\,
            in2 => \_gnd_net_\,
            in3 => \N__23510\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__47779\,
            ce => 'H',
            sr => \N__47416\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26958\,
            in1 => \N__25223\,
            in2 => \_gnd_net_\,
            in3 => \N__23507\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47779\,
            ce => 'H',
            sr => \N__47416\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26225\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25687\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25378\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25546\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25888\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26121\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33377\,
            in2 => \_gnd_net_\,
            in3 => \N__33851\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_434_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30514\,
            in2 => \N__30518\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__27975\,
            in1 => \N__25615\,
            in2 => \N__25592\,
            in3 => \N__23540\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            clk => \N__47852\,
            ce => 'H',
            sr => \N__47327\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__27965\,
            in1 => \N__30527\,
            in2 => \N__28370\,
            in3 => \N__23537\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            clk => \N__47852\,
            ce => 'H',
            sr => \N__47327\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__27976\,
            in1 => \N__26138\,
            in2 => \N__25574\,
            in3 => \N__23534\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            clk => \N__47852\,
            ce => 'H',
            sr => \N__47327\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0111110111010111"
        )
    port map (
            in0 => \N__27966\,
            in1 => \N__23531\,
            in2 => \N__25394\,
            in3 => \N__23525\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            clk => \N__47852\,
            ce => 'H',
            sr => \N__47327\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25178\,
            in2 => \N__25457\,
            in3 => \N__23522\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23744\,
            in2 => \N__23738\,
            in3 => \N__23717\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23714\,
            in2 => \N__28382\,
            in3 => \N__23693\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23690\,
            in2 => \N__23684\,
            in3 => \N__23666\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30728\,
            in2 => \N__25583\,
            in3 => \N__23663\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23660\,
            in2 => \N__25916\,
            in3 => \N__23639\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23636\,
            in2 => \N__25970\,
            in3 => \N__23615\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23612\,
            in2 => \N__25466\,
            in3 => \N__23600\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25517\,
            in2 => \N__28442\,
            in3 => \N__23597\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40502\,
            in2 => \N__25961\,
            in3 => \N__23861\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23858\,
            in2 => \N__25526\,
            in3 => \N__23849\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24002\,
            in2 => \N__24059\,
            in3 => \N__23837\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23834\,
            in2 => \N__25334\,
            in3 => \N__23819\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23816\,
            in2 => \N__25817\,
            in3 => \N__23798\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23795\,
            in2 => \N__25865\,
            in3 => \N__23777\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28505\,
            in2 => \N__26246\,
            in3 => \N__23768\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23765\,
            in2 => \N__26189\,
            in3 => \N__23747\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30653\,
            in2 => \N__25805\,
            in3 => \N__23972\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23993\,
            in2 => \N__26027\,
            in3 => \N__23960\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23957\,
            in2 => \N__26327\,
            in3 => \N__23939\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30449\,
            in2 => \N__26315\,
            in3 => \N__23930\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26258\,
            in2 => \N__25628\,
            in3 => \N__23918\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26078\,
            in2 => \N__23915\,
            in3 => \N__23897\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23894\,
            in2 => \N__29231\,
            in3 => \N__23873\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24065\,
            in2 => \N__33503\,
            in3 => \N__23864\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33501\,
            in2 => \N__24107\,
            in3 => \N__24161\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33502\,
            in2 => \N__40565\,
            in3 => \N__24152\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28233\,
            in1 => \N__33727\,
            in2 => \_gnd_net_\,
            in3 => \N__24149\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24126\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24084\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29013\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33725\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24045\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__24046\,
            in1 => \N__33726\,
            in2 => \N__28897\,
            in3 => \N__28871\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26061\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33743\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29108\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28896\,
            in2 => \_gnd_net_\,
            in3 => \N__33742\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36301\,
            in2 => \_gnd_net_\,
            in3 => \N__36254\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__24449\,
            in1 => \N__27122\,
            in2 => \N__35816\,
            in3 => \N__24482\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__24336\,
            sr => \N__47365\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27339\,
            in1 => \N__27114\,
            in2 => \N__27505\,
            in3 => \N__24450\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__24336\,
            sr => \N__47365\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__27111\,
            in1 => \N__26617\,
            in2 => \_gnd_net_\,
            in3 => \N__27342\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__24336\,
            sr => \N__47365\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__27337\,
            in1 => \N__26647\,
            in2 => \_gnd_net_\,
            in3 => \N__27115\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__24336\,
            sr => \N__47365\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__27110\,
            in1 => \N__27340\,
            in2 => \_gnd_net_\,
            in3 => \N__26675\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__24336\,
            sr => \N__47365\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__27336\,
            in1 => \N__27113\,
            in2 => \_gnd_net_\,
            in3 => \N__33939\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__24336\,
            sr => \N__47365\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__27112\,
            in1 => \N__27341\,
            in2 => \N__27836\,
            in3 => \N__27196\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__24336\,
            sr => \N__47365\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27338\,
            in1 => \N__26864\,
            in2 => \_gnd_net_\,
            in3 => \N__24945\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__24336\,
            sr => \N__47365\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26429\,
            in2 => \_gnd_net_\,
            in3 => \N__26749\,
            lcout => \elapsed_time_ns_1_RNI62CED1_0_19\,
            ltout => \elapsed_time_ns_1_RNI62CED1_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27355\,
            in2 => \N__24254\,
            in3 => \N__27118\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47804\,
            ce => \N__27023\,
            sr => \N__47374\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__27832\,
            in1 => \N__27426\,
            in2 => \_gnd_net_\,
            in3 => \N__27188\,
            lcout => \phase_controller_inst1.stoper_hc.N_315\,
            ltout => \phase_controller_inst1.stoper_hc.N_315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__31246\,
            in1 => \N__27356\,
            in2 => \N__24251\,
            in3 => \N__27119\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47804\,
            ce => \N__27023\,
            sr => \N__47374\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24459\,
            in1 => \N__27357\,
            in2 => \N__27469\,
            in3 => \N__27117\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47804\,
            ce => \N__27023\,
            sr => \N__47374\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27116\,
            in1 => \N__27358\,
            in2 => \N__24467\,
            in3 => \N__27509\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47804\,
            ce => \N__27023\,
            sr => \N__47374\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__35927\,
            in1 => \N__26648\,
            in2 => \N__31958\,
            in3 => \N__36974\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24248\,
            in3 => \N__26752\,
            lcout => \elapsed_time_ns_1_RNI51CED1_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__27251\,
            in1 => \N__37147\,
            in2 => \N__36996\,
            in3 => \N__31791\,
            lcout => \elapsed_time_ns_1_RNIQ4OD11_0_31\,
            ltout => \elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1_9_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110010"
        )
    port map (
            in0 => \N__27365\,
            in1 => \N__27105\,
            in2 => \N__24485\,
            in3 => \N__26591\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__35815\,
            in1 => \N__27121\,
            in2 => \N__24473\,
            in3 => \N__24458\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__27022\,
            sr => \N__47380\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__27427\,
            in1 => \N__27106\,
            in2 => \N__24468\,
            in3 => \N__27255\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__27022\,
            sr => \N__47380\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__27529\,
            in1 => \N__27120\,
            in2 => \N__27299\,
            in3 => \N__24457\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__27022\,
            sr => \N__47380\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__27266\,
            in1 => \N__24557\,
            in2 => \N__26576\,
            in3 => \N__27148\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001111"
        )
    port map (
            in0 => \N__26537\,
            in1 => \N__24555\,
            in2 => \N__37256\,
            in3 => \N__26574\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26536\,
            in2 => \_gnd_net_\,
            in3 => \N__37252\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.N_283_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27147\,
            in1 => \N__24556\,
            in2 => \N__24392\,
            in3 => \N__26575\,
            lcout => \phase_controller_inst1.stoper_hc.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__35926\,
            in1 => \N__24576\,
            in2 => \N__31871\,
            in3 => \N__36970\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24584\,
            in3 => \N__26751\,
            lcout => \elapsed_time_ns_1_RNIIU2KD1_0_6\,
            ltout => \elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__27376\,
            in1 => \N__26819\,
            in2 => \N__24560\,
            in3 => \N__26847\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__27146\,
            in1 => \_gnd_net_\,
            in2 => \N__24542\,
            in3 => \N__27819\,
            lcout => \phase_controller_inst1.stoper_hc.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001110"
        )
    port map (
            in0 => \N__27192\,
            in1 => \N__27383\,
            in2 => \N__27160\,
            in3 => \N__27818\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24515\,
            in2 => \N__24539\,
            in3 => \N__27300\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111101110"
        )
    port map (
            in0 => \N__24516\,
            in1 => \N__35928\,
            in2 => \N__31574\,
            in3 => \N__37001\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24521\,
            in3 => \N__26756\,
            lcout => \elapsed_time_ns_1_RNIDP2KD1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__24861\,
            in1 => \N__24496\,
            in2 => \N__24949\,
            in3 => \N__27304\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47789\,
            ce => \N__27014\,
            sr => \N__47393\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__26698\,
            in1 => \N__24925\,
            in2 => \N__27343\,
            in3 => \N__24862\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47789\,
            ce => \N__27014\,
            sr => \N__47393\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24818\,
            in2 => \N__24779\,
            in3 => \N__24806\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24770\,
            in2 => \N__24752\,
            in3 => \N__24763\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24742\,
            in1 => \N__24731\,
            in2 => \N__24719\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24710\,
            in1 => \N__24692\,
            in2 => \N__24686\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24674\,
            in2 => \N__24653\,
            in3 => \N__24664\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24643\,
            in1 => \N__24620\,
            in2 => \N__24632\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24590\,
            in2 => \N__24614\,
            in3 => \N__24601\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25145\,
            in2 => \N__25172\,
            in3 => \N__25160\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25115\,
            in2 => \N__25139\,
            in3 => \N__25126\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25109\,
            in2 => \N__25088\,
            in3 => \N__25099\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25079\,
            in2 => \N__25055\,
            in3 => \N__25066\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25022\,
            in2 => \N__25046\,
            in3 => \N__25033\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25016\,
            in2 => \N__24995\,
            in3 => \N__25006\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24983\,
            in2 => \N__24962\,
            in3 => \N__24973\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25324\,
            in1 => \N__25313\,
            in2 => \N__27035\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25307\,
            in2 => \N__25286\,
            in3 => \N__25297\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26462\,
            in2 => \N__25265\,
            in3 => \N__25276\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25256\,
            in2 => \N__25232\,
            in3 => \N__25243\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25222\,
            in1 => \N__25199\,
            in2 => \N__25211\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25193\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32418\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47767\,
            ce => 'H',
            sr => \N__47418\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__25736\,
            in1 => \N__31090\,
            in2 => \N__33775\,
            in3 => \N__28760\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25735\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__28308\,
            in1 => \N__28158\,
            in2 => \N__27999\,
            in3 => \N__25445\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => 'H',
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__28156\,
            in1 => \N__28309\,
            in2 => \N__25439\,
            in3 => \N__27974\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => 'H',
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__27967\,
            in1 => \N__25430\,
            in2 => \N__28319\,
            in3 => \N__28159\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => 'H',
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25548\,
            in1 => \N__40519\,
            in2 => \N__28479\,
            in3 => \N__28306\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__28307\,
            in1 => \N__28157\,
            in2 => \N__27998\,
            in3 => \N__25412\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => 'H',
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25547\,
            in1 => \N__40520\,
            in2 => \N__28478\,
            in3 => \N__40605\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__25697\,
            in1 => \N__33695\,
            in2 => \N__30830\,
            in3 => \N__28769\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__25382\,
            in1 => \N__30644\,
            in2 => \N__33757\,
            in3 => \N__28859\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26298\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33692\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28636\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__25616\,
            in1 => \N__33693\,
            in2 => \N__30923\,
            in3 => \N__28538\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__30767\,
            in1 => \N__28696\,
            in2 => \N__33756\,
            in3 => \N__28679\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__26165\,
            in1 => \N__33694\,
            in2 => \N__30868\,
            in3 => \N__28514\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__28937\,
            in1 => \N__25558\,
            in2 => \N__28913\,
            in3 => \N__33712\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__28483\,
            in1 => \N__28991\,
            in2 => \N__33759\,
            in3 => \N__29015\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29036\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33703\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__33708\,
            in1 => \N__25505\,
            in2 => \N__25469\,
            in3 => \N__29024\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__28635\,
            in1 => \N__26013\,
            in2 => \N__28616\,
            in3 => \N__33707\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011111111"
        )
    port map (
            in0 => \N__40536\,
            in1 => \N__28979\,
            in2 => \N__28952\,
            in3 => \N__33741\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28697\,
            in2 => \_gnd_net_\,
            in3 => \N__33702\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__25952\,
            in1 => \N__28663\,
            in2 => \N__33758\,
            in3 => \N__28646\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__25906\,
            in1 => \N__33718\,
            in2 => \N__28808\,
            in3 => \N__28778\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33760\,
            in3 => \N__28667\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__25856\,
            in1 => \N__33717\,
            in2 => \N__28847\,
            in3 => \N__28817\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__31361\,
            in1 => \N__30698\,
            in2 => \N__33761\,
            in3 => \N__29132\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__25796\,
            in1 => \N__25746\,
            in2 => \N__25715\,
            in3 => \N__25664\,
            lcout => \current_shift_inst.PI_CTRL.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33716\,
            in1 => \N__29165\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__33755\,
            in1 => \N__27598\,
            in2 => \N__26249\,
            in3 => \N__29153\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111101101111"
        )
    port map (
            in0 => \N__31289\,
            in1 => \N__29144\,
            in2 => \N__33762\,
            in3 => \N__26236\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__28933\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33669\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26175\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29057\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33670\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__33676\,
            in1 => \N__26125\,
            in2 => \N__26081\,
            in3 => \N__29045\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__31313\,
            in1 => \N__26071\,
            in2 => \N__29120\,
            in3 => \N__33671\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__26506\,
            in1 => \N__37154\,
            in2 => \N__31703\,
            in3 => \N__36981\,
            lcout => \elapsed_time_ns_1_RNIP2ND11_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__29106\,
            in1 => \N__26366\,
            in2 => \N__29087\,
            in3 => \N__33672\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__30499\,
            in1 => \N__31388\,
            in2 => \N__33745\,
            in3 => \N__29075\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__31793\,
            in1 => \N__31526\,
            in2 => \N__31844\,
            in3 => \N__31817\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__31898\,
            in1 => \N__27404\,
            in2 => \N__26306\,
            in3 => \N__36897\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26303\,
            in3 => \N__26735\,
            lcout => \elapsed_time_ns_1_RNI1TBED1_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__37102\,
            in1 => \N__26393\,
            in2 => \N__29402\,
            in3 => \N__36895\,
            lcout => \elapsed_time_ns_1_RNIV8ND11_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101101111011"
        )
    port map (
            in0 => \N__29066\,
            in1 => \N__33744\,
            in2 => \N__31337\,
            in3 => \N__26299\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__37103\,
            in1 => \N__26378\,
            in2 => \N__29426\,
            in3 => \N__36896\,
            lcout => \elapsed_time_ns_1_RNIU7ND11_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26734\,
            in2 => \_gnd_net_\,
            in3 => \N__35780\,
            lcout => \elapsed_time_ns_1_RNIL13KD1_0_9\,
            ltout => \elapsed_time_ns_1_RNIL13KD1_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_9_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27831\,
            in2 => \N__26423\,
            in3 => \N__27403\,
            lcout => \phase_controller_inst1.stoper_hc.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__37075\,
            in1 => \N__26420\,
            in2 => \N__29348\,
            in3 => \N__36864\,
            lcout => \elapsed_time_ns_1_RNI1BND11_0_29\,
            ltout => \elapsed_time_ns_1_RNI1BND11_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26414\,
            in3 => \N__29212\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__47479\,
            in1 => \N__29171\,
            in2 => \N__31792\,
            in3 => \N__29195\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__36867\,
            in1 => \N__37078\,
            in2 => \N__31445\,
            in3 => \N__27503\,
            lcout => \elapsed_time_ns_1_RNIQ2MD11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__37077\,
            in1 => \N__26402\,
            in2 => \N__29375\,
            in3 => \N__36866\,
            lcout => \elapsed_time_ns_1_RNI0AND11_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__36868\,
            in1 => \N__26492\,
            in2 => \N__37153\,
            in3 => \N__29468\,
            lcout => \elapsed_time_ns_1_RNIS5ND11_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__37076\,
            in1 => \N__36865\,
            in2 => \N__26411\,
            in3 => \N__29450\,
            lcout => \elapsed_time_ns_1_RNIT6ND11_0_25\,
            ltout => \elapsed_time_ns_1_RNIT6ND11_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26401\,
            in1 => \N__26392\,
            in2 => \N__26381\,
            in3 => \N__26377\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26437\,
            in1 => \N__26449\,
            in2 => \N__26510\,
            in3 => \N__26491\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26480\,
            in1 => \N__36815\,
            in2 => \N__26474\,
            in3 => \N__26471\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27298\,
            in2 => \N__26465\,
            in3 => \N__26673\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47795\,
            ce => \N__27013\,
            sr => \N__47358\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__26450\,
            in1 => \N__37106\,
            in2 => \N__31721\,
            in3 => \N__36898\,
            lcout => \elapsed_time_ns_1_RNIQ3ND11_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__26674\,
            in1 => \N__36899\,
            in2 => \N__35922\,
            in3 => \N__31973\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26441\,
            in3 => \N__26748\,
            lcout => \elapsed_time_ns_1_RNI40CED1_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__37105\,
            in1 => \N__26438\,
            in2 => \N__36994\,
            in3 => \N__29486\,
            lcout => \elapsed_time_ns_1_RNIR4ND11_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010111010"
        )
    port map (
            in0 => \N__35918\,
            in1 => \N__36969\,
            in2 => \N__26618\,
            in3 => \N__31926\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35917\,
            in2 => \_gnd_net_\,
            in3 => \N__26516\,
            lcout => \elapsed_time_ns_1_RNIQURR91_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26561\,
            in1 => \N__27545\,
            in2 => \N__29446\,
            in3 => \N__29464\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33878\,
            in2 => \_gnd_net_\,
            in3 => \N__26750\,
            lcout => \elapsed_time_ns_1_RNI3VBED1_0_16\,
            ltout => \elapsed_time_ns_1_RNI3VBED1_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__26671\,
            in1 => \N__26638\,
            in2 => \N__26705\,
            in3 => \N__26612\,
            lcout => \phase_controller_inst1.stoper_hc.N_278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__37146\,
            in1 => \N__31592\,
            in2 => \N__36995\,
            in3 => \N__26691\,
            lcout => \elapsed_time_ns_1_RNIA3DJ11_0_4\,
            ltout => \elapsed_time_ns_1_RNIA3DJ11_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26672\,
            in1 => \N__26787\,
            in2 => \N__26651\,
            in3 => \N__33929\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__26639\,
            in1 => \N__26613\,
            in2 => \N__26594\,
            in3 => \N__26590\,
            lcout => \phase_controller_inst1.stoper_hc.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111110"
        )
    port map (
            in0 => \N__29416\,
            in1 => \N__29389\,
            in2 => \N__29368\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__36961\,
            in1 => \N__37145\,
            in2 => \N__31499\,
            in3 => \N__27448\,
            lcout => \elapsed_time_ns_1_RNIP1MD11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__31547\,
            in1 => \N__31985\,
            in2 => \N__26555\,
            in3 => \N__36962\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29338\,
            in1 => \N__29482\,
            in2 => \N__37018\,
            in3 => \N__29653\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__27525\,
            in1 => \N__31484\,
            in2 => \N__36982\,
            in3 => \N__37144\,
            lcout => \elapsed_time_ns_1_RNINVLD11_0_10\,
            ltout => \elapsed_time_ns_1_RNINVLD11_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31245\,
            in1 => \N__27504\,
            in2 => \N__27473\,
            in3 => \N__27447\,
            lcout => \phase_controller_inst1.stoper_hc.N_319\,
            ltout => \phase_controller_inst1.stoper_hc.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111111"
        )
    port map (
            in0 => \N__35820\,
            in1 => \_gnd_net_\,
            in2 => \N__27434\,
            in3 => \N__27416\,
            lcout => \phase_controller_inst1.stoper_hc.N_275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0_9_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__27817\,
            in1 => \N__35821\,
            in2 => \_gnd_net_\,
            in3 => \N__27377\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a5_1_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__27820\,
            in1 => \N__27305\,
            in2 => \N__27197\,
            in3 => \N__27142\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47781\,
            ce => \N__27016\,
            sr => \N__47381\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__37143\,
            in1 => \N__31166\,
            in2 => \N__37000\,
            in3 => \N__26853\,
            lcout => \elapsed_time_ns_1_RNID6DJ11_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__37142\,
            in1 => \N__31187\,
            in2 => \N__36999\,
            in3 => \N__26826\,
            lcout => \elapsed_time_ns_1_RNIE7DJ11_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__37141\,
            in1 => \N__36984\,
            in2 => \N__31613\,
            in3 => \N__26786\,
            lcout => \elapsed_time_ns_1_RNIB4DJ11_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__31211\,
            in1 => \N__27821\,
            in2 => \N__37155\,
            in3 => \N__36983\,
            lcout => \elapsed_time_ns_1_RNIS4MD11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNI8HMG_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27706\,
            in1 => \N__27751\,
            in2 => \_gnd_net_\,
            in3 => \N__27781\,
            lcout => \phase_controller_inst2.stoper_hc.running_1_sqmuxa\,
            ltout => \phase_controller_inst2.stoper_hc.running_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__27752\,
            in1 => \N__27707\,
            in2 => \N__27674\,
            in3 => \N__27671\,
            lcout => \phase_controller_inst2.stoper_hc.un1_start_latched2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34043\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47761\,
            ce => 'H',
            sr => \N__47417\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27629\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27605\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28800\,
            in2 => \_gnd_net_\,
            in3 => \N__33763\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27595\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28465\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__28427\,
            in1 => \N__31024\,
            in2 => \N__28727\,
            in3 => \N__33765\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__33764\,
            in1 => \N__30558\,
            in2 => \N__28529\,
            in3 => \N__30892\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36161\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__47318\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28574\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__47318\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30829\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__47318\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30983\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__47318\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__28328\,
            in1 => \N__28318\,
            in2 => \N__28166\,
            in3 => \N__27997\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__47318\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30922\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__47318\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30893\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__47318\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28562\,
            in2 => \_gnd_net_\,
            in3 => \N__28573\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30979\,
            in1 => \N__28556\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28550\,
            in2 => \_gnd_net_\,
            in3 => \N__30961\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28544\,
            in2 => \_gnd_net_\,
            in3 => \N__30937\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30995\,
            in2 => \_gnd_net_\,
            in3 => \N__28532\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30716\,
            in2 => \_gnd_net_\,
            in3 => \N__28517\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30704\,
            in2 => \_gnd_net_\,
            in3 => \N__28508\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30788\,
            in2 => \_gnd_net_\,
            in3 => \N__28763\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31067\,
            in2 => \_gnd_net_\,
            in3 => \N__28745\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_8\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31034\,
            in2 => \_gnd_net_\,
            in3 => \N__28730\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31001\,
            in2 => \_gnd_net_\,
            in3 => \N__28715\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30710\,
            in2 => \_gnd_net_\,
            in3 => \N__28700\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28695\,
            in2 => \_gnd_net_\,
            in3 => \N__28670\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28662\,
            in2 => \_gnd_net_\,
            in3 => \N__28640\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28637\,
            in2 => \_gnd_net_\,
            in3 => \N__28607\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29035\,
            in2 => \_gnd_net_\,
            in3 => \N__29018\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29014\,
            in2 => \_gnd_net_\,
            in3 => \N__28982\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28975\,
            in2 => \_gnd_net_\,
            in3 => \N__28940\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28929\,
            in2 => \_gnd_net_\,
            in3 => \N__28901\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28898\,
            in2 => \_gnd_net_\,
            in3 => \N__28862\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30640\,
            in2 => \_gnd_net_\,
            in3 => \N__28850\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28840\,
            in2 => \_gnd_net_\,
            in3 => \N__28811\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28801\,
            in2 => \_gnd_net_\,
            in3 => \N__28772\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29164\,
            in2 => \_gnd_net_\,
            in3 => \N__29147\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31281\,
            in2 => \_gnd_net_\,
            in3 => \N__29135\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31353\,
            in2 => \_gnd_net_\,
            in3 => \N__29123\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31305\,
            in2 => \_gnd_net_\,
            in3 => \N__29111\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29107\,
            in2 => \_gnd_net_\,
            in3 => \N__29078\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31384\,
            in3 => \N__29069\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31329\,
            in2 => \_gnd_net_\,
            in3 => \N__29060\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29056\,
            in2 => \_gnd_net_\,
            in3 => \N__29039\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__29273\,
            in1 => \N__33602\,
            in2 => \_gnd_net_\,
            in3 => \N__29234\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__32003\,
            in1 => \N__47476\,
            in2 => \N__31622\,
            in3 => \N__31505\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__32002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31732\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_382_i\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_382_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__29213\,
            in1 => \N__29660\,
            in2 => \N__29216\,
            in3 => \N__37131\,
            lcout => \elapsed_time_ns_1_RNIP3OD11_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__35845\,
            in1 => \N__31183\,
            in2 => \_gnd_net_\,
            in3 => \N__31162\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__31894\,
            in1 => \N__31210\,
            in2 => \N__29201\,
            in3 => \N__31423\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110011"
        )
    port map (
            in0 => \N__31904\,
            in1 => \N__31681\,
            in2 => \N__29198\,
            in3 => \N__29188\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__31682\,
            in1 => \N__47475\,
            in2 => \N__29189\,
            in3 => \N__32001\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__31519\,
            in1 => \N__29184\,
            in2 => \_gnd_net_\,
            in3 => \N__31403\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29636\,
            in2 => \N__29608\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47790\,
            ce => \N__37177\,
            sr => \N__47349\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37225\,
            in2 => \N__29576\,
            in3 => \N__29297\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47790\,
            ce => \N__37177\,
            sr => \N__47349\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29609\,
            in2 => \N__29545\,
            in3 => \N__29294\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47790\,
            ce => \N__37177\,
            sr => \N__47349\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29575\,
            in2 => \N__29518\,
            in3 => \N__29291\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47790\,
            ce => \N__37177\,
            sr => \N__47349\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29884\,
            in2 => \N__29546\,
            in3 => \N__29288\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47790\,
            ce => \N__37177\,
            sr => \N__47349\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29857\,
            in2 => \N__29519\,
            in3 => \N__29285\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47790\,
            ce => \N__37177\,
            sr => \N__47349\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29827\,
            in2 => \N__29888\,
            in3 => \N__29282\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47790\,
            ce => \N__37177\,
            sr => \N__47349\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29858\,
            in2 => \N__29800\,
            in3 => \N__29279\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47790\,
            ce => \N__37177\,
            sr => \N__47349\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29767\,
            in2 => \N__29834\,
            in3 => \N__29276\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47785\,
            ce => \N__37176\,
            sr => \N__47359\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29801\,
            in2 => \N__29743\,
            in3 => \N__29324\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47785\,
            ce => \N__37176\,
            sr => \N__47359\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29768\,
            in2 => \N__29716\,
            in3 => \N__29321\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47785\,
            ce => \N__37176\,
            sr => \N__47359\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29686\,
            in2 => \N__29744\,
            in3 => \N__29318\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47785\,
            ce => \N__37176\,
            sr => \N__47359\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30106\,
            in2 => \N__29717\,
            in3 => \N__29315\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47785\,
            ce => \N__37176\,
            sr => \N__47359\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30079\,
            in2 => \N__29690\,
            in3 => \N__29312\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47785\,
            ce => \N__37176\,
            sr => \N__47359\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30052\,
            in2 => \N__30110\,
            in3 => \N__29309\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47785\,
            ce => \N__37176\,
            sr => \N__47359\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30080\,
            in2 => \N__30022\,
            in3 => \N__29306\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47785\,
            ce => \N__37176\,
            sr => \N__47359\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29986\,
            in2 => \N__30056\,
            in3 => \N__29303\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47782\,
            ce => \N__37175\,
            sr => \N__47366\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29959\,
            in2 => \N__30023\,
            in3 => \N__29300\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47782\,
            ce => \N__37175\,
            sr => \N__47366\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29938\,
            in2 => \N__29990\,
            in3 => \N__29492\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47782\,
            ce => \N__37175\,
            sr => \N__47366\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29960\,
            in2 => \N__29918\,
            in3 => \N__29489\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47782\,
            ce => \N__37175\,
            sr => \N__47366\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29939\,
            in2 => \N__30436\,
            in3 => \N__29471\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47782\,
            ce => \N__37175\,
            sr => \N__47366\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29917\,
            in2 => \N__30409\,
            in3 => \N__29453\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47782\,
            ce => \N__37175\,
            sr => \N__47366\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30379\,
            in2 => \N__30437\,
            in3 => \N__29429\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47782\,
            ce => \N__37175\,
            sr => \N__47366\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30355\,
            in2 => \N__30410\,
            in3 => \N__29405\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47782\,
            ce => \N__37175\,
            sr => \N__47366\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30325\,
            in2 => \N__30383\,
            in3 => \N__29378\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47777\,
            ce => \N__37174\,
            sr => \N__47375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30356\,
            in2 => \N__30298\,
            in3 => \N__29351\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47777\,
            ce => \N__37174\,
            sr => \N__47375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30272\,
            in2 => \N__30329\,
            in3 => \N__29327\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47777\,
            ce => \N__37174\,
            sr => \N__47375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30251\,
            in2 => \N__30299\,
            in3 => \N__29642\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47777\,
            ce => \N__37174\,
            sr => \N__47375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29639\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47777\,
            ce => \N__37174\,
            sr => \N__47375\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29635\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47777\,
            ce => \N__37174\,
            sr => \N__47375\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30233\,
            in1 => \N__29631\,
            in2 => \_gnd_net_\,
            in3 => \N__29615\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__47772\,
            ce => \N__32312\,
            sr => \N__47382\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30229\,
            in1 => \N__37218\,
            in2 => \_gnd_net_\,
            in3 => \N__29612\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__47772\,
            ce => \N__32312\,
            sr => \N__47382\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30234\,
            in1 => \N__29601\,
            in2 => \_gnd_net_\,
            in3 => \N__29579\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__47772\,
            ce => \N__32312\,
            sr => \N__47382\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30230\,
            in1 => \N__29565\,
            in2 => \_gnd_net_\,
            in3 => \N__29549\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__47772\,
            ce => \N__32312\,
            sr => \N__47382\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30235\,
            in1 => \N__29538\,
            in2 => \_gnd_net_\,
            in3 => \N__29522\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__47772\,
            ce => \N__32312\,
            sr => \N__47382\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30231\,
            in1 => \N__29506\,
            in2 => \_gnd_net_\,
            in3 => \N__29891\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__47772\,
            ce => \N__32312\,
            sr => \N__47382\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30236\,
            in1 => \N__29877\,
            in2 => \_gnd_net_\,
            in3 => \N__29861\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__47772\,
            ce => \N__32312\,
            sr => \N__47382\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30232\,
            in1 => \N__29851\,
            in2 => \_gnd_net_\,
            in3 => \N__29837\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__47772\,
            ce => \N__32312\,
            sr => \N__47382\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30220\,
            in1 => \N__29826\,
            in2 => \_gnd_net_\,
            in3 => \N__29804\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__47769\,
            ce => \N__32307\,
            sr => \N__47388\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30224\,
            in1 => \N__29793\,
            in2 => \_gnd_net_\,
            in3 => \N__29771\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__47769\,
            ce => \N__32307\,
            sr => \N__47388\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30217\,
            in1 => \N__29761\,
            in2 => \_gnd_net_\,
            in3 => \N__29747\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__47769\,
            ce => \N__32307\,
            sr => \N__47388\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30221\,
            in1 => \N__29736\,
            in2 => \_gnd_net_\,
            in3 => \N__29720\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__47769\,
            ce => \N__32307\,
            sr => \N__47388\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30218\,
            in1 => \N__29709\,
            in2 => \_gnd_net_\,
            in3 => \N__29693\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__47769\,
            ce => \N__32307\,
            sr => \N__47388\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30222\,
            in1 => \N__29679\,
            in2 => \_gnd_net_\,
            in3 => \N__29663\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__47769\,
            ce => \N__32307\,
            sr => \N__47388\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30219\,
            in1 => \N__30099\,
            in2 => \_gnd_net_\,
            in3 => \N__30083\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__47769\,
            ce => \N__32307\,
            sr => \N__47388\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30223\,
            in1 => \N__30073\,
            in2 => \_gnd_net_\,
            in3 => \N__30059\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__47769\,
            ce => \N__32307\,
            sr => \N__47388\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30213\,
            in1 => \N__30045\,
            in2 => \_gnd_net_\,
            in3 => \N__30026\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__47764\,
            ce => \N__32311\,
            sr => \N__47394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30225\,
            in1 => \N__30009\,
            in2 => \_gnd_net_\,
            in3 => \N__29993\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__47764\,
            ce => \N__32311\,
            sr => \N__47394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30214\,
            in1 => \N__29979\,
            in2 => \_gnd_net_\,
            in3 => \N__29963\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__47764\,
            ce => \N__32311\,
            sr => \N__47394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30226\,
            in1 => \N__29958\,
            in2 => \_gnd_net_\,
            in3 => \N__29942\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__47764\,
            ce => \N__32311\,
            sr => \N__47394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30215\,
            in1 => \N__29937\,
            in2 => \_gnd_net_\,
            in3 => \N__29921\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__47764\,
            ce => \N__32311\,
            sr => \N__47394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30227\,
            in1 => \N__29913\,
            in2 => \_gnd_net_\,
            in3 => \N__29894\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__47764\,
            ce => \N__32311\,
            sr => \N__47394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30216\,
            in1 => \N__30429\,
            in2 => \_gnd_net_\,
            in3 => \N__30413\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__47764\,
            ce => \N__32311\,
            sr => \N__47394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30228\,
            in1 => \N__30402\,
            in2 => \_gnd_net_\,
            in3 => \N__30386\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__47764\,
            ce => \N__32311\,
            sr => \N__47394\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30189\,
            in1 => \N__30378\,
            in2 => \_gnd_net_\,
            in3 => \N__30359\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__47762\,
            ce => \N__32294\,
            sr => \N__47399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30193\,
            in1 => \N__30348\,
            in2 => \_gnd_net_\,
            in3 => \N__30332\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__47762\,
            ce => \N__32294\,
            sr => \N__47399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30190\,
            in1 => \N__30318\,
            in2 => \_gnd_net_\,
            in3 => \N__30302\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__47762\,
            ce => \N__32294\,
            sr => \N__47399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30194\,
            in1 => \N__30291\,
            in2 => \_gnd_net_\,
            in3 => \N__30275\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__47762\,
            ce => \N__32294\,
            sr => \N__47399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30191\,
            in1 => \N__30271\,
            in2 => \_gnd_net_\,
            in3 => \N__30257\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__47762\,
            ce => \N__32294\,
            sr => \N__47399\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__30250\,
            in1 => \N__30192\,
            in2 => \_gnd_net_\,
            in3 => \N__30254\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47762\,
            ce => \N__32294\,
            sr => \N__47399\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32217\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32216\,
            in2 => \_gnd_net_\,
            in3 => \N__32246\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_432_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30587\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30599\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32267\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30580\,
            ce => 'H',
            sr => \N__47299\
        );

    \delay_measurement_inst.stop_timer_hc_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32268\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30581\,
            ce => 'H',
            sr => \N__47304\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30557\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33766\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30495\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33376\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30965\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47817\,
            ce => 'H',
            sr => \N__47314\
        );

    \phase_controller_inst1.stoper_tr.running_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000101110"
        )
    port map (
            in0 => \N__42900\,
            in1 => \N__42845\,
            in2 => \N__42980\,
            in3 => \N__43043\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47817\,
            ce => 'H',
            sr => \N__47314\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30814\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30746\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30885\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31119\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30849\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30696\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__30639\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33679\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30907\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30989\,
            in2 => \_gnd_net_\,
            in3 => \N__36157\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35942\,
            in2 => \_gnd_net_\,
            in3 => \N__30968\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__47805\,
            ce => 'H',
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31265\,
            in2 => \_gnd_net_\,
            in3 => \N__30950\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__47805\,
            ce => 'H',
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31397\,
            in2 => \_gnd_net_\,
            in3 => \N__30926\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__47805\,
            ce => 'H',
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33956\,
            in3 => \N__30896\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__47805\,
            ce => 'H',
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34523\,
            in2 => \_gnd_net_\,
            in3 => \N__30872\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__47805\,
            ce => 'H',
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33788\,
            in2 => \_gnd_net_\,
            in3 => \N__30833\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__47805\,
            ce => 'H',
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34571\,
            in2 => \_gnd_net_\,
            in3 => \N__31145\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__47805\,
            ce => 'H',
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33293\,
            in2 => \_gnd_net_\,
            in3 => \N__31142\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__47801\,
            ce => 'H',
            sr => \N__47328\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33476\,
            in2 => \_gnd_net_\,
            in3 => \N__31139\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__47801\,
            ce => 'H',
            sr => \N__47328\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32324\,
            in2 => \_gnd_net_\,
            in3 => \N__31136\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__47801\,
            ce => 'H',
            sr => \N__47328\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33863\,
            in2 => \_gnd_net_\,
            in3 => \N__31100\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__47801\,
            ce => 'H',
            sr => \N__47328\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36671\,
            in2 => \_gnd_net_\,
            in3 => \N__31097\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47801\,
            ce => 'H',
            sr => \N__47328\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31078\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31045\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31012\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36512\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31383\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33600\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33598\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31357\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31333\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33601\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33599\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31309\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31285\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33597\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36125\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__31235\,
            in1 => \N__36934\,
            in2 => \N__31469\,
            in3 => \N__37104\,
            lcout => \elapsed_time_ns_1_RNIO0MD11_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31209\,
            in1 => \N__31182\,
            in2 => \N__31427\,
            in3 => \N__31161\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__35844\,
            in1 => \N__31580\,
            in2 => \N__31631\,
            in3 => \N__31628\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__31539\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37201\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47474\,
            in1 => \N__31786\,
            in2 => \_gnd_net_\,
            in3 => \N__31813\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31603\,
            in2 => \_gnd_net_\,
            in3 => \N__31591\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37202\,
            in1 => \N__31573\,
            in2 => \N__31550\,
            in3 => \N__31540\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__31787\,
            in1 => \N__47473\,
            in2 => \N__31508\,
            in3 => \N__31837\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31495\,
            in1 => \N__31480\,
            in2 => \N__31462\,
            in3 => \N__31438\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__47477\,
            in1 => \N__31833\,
            in2 => \N__31675\,
            in3 => \N__31409\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31887\,
            in1 => \N__31861\,
            in2 => \N__33898\,
            in3 => \N__31951\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31972\,
            in1 => \N__31934\,
            in2 => \N__32012\,
            in3 => \N__32009\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__31733\,
            in1 => \_gnd_net_\,
            in2 => \N__31988\,
            in3 => \N__47478\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31971\,
            in1 => \N__31950\,
            in2 => \N__31933\,
            in3 => \N__33891\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31886\,
            in1 => \N__31860\,
            in2 => \N__31847\,
            in3 => \N__35843\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__31812\,
            in1 => \_gnd_net_\,
            in2 => \N__31796\,
            in3 => \N__31771\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31714\,
            in2 => \_gnd_net_\,
            in3 => \N__31693\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__33847\,
            in1 => \N__33360\,
            in2 => \_gnd_net_\,
            in3 => \N__33821\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => 'H',
            sr => \N__47350\
        );

    \phase_controller_inst2.T01_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__31642\,
            in1 => \N__32398\,
            in2 => \_gnd_net_\,
            in3 => \N__32148\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => 'H',
            sr => \N__47350\
        );

    \phase_controller_inst2.T12_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__32167\,
            in1 => \N__34029\,
            in2 => \_gnd_net_\,
            in3 => \N__32149\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => 'H',
            sr => \N__47350\
        );

    \phase_controller_inst2.state_1_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__33996\,
            in1 => \N__32156\,
            in2 => \N__32123\,
            in3 => \N__34027\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => 'H',
            sr => \N__47360\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34696\,
            in2 => \_gnd_net_\,
            in3 => \N__34656\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__32362\,
            in1 => \N__34028\,
            in2 => \N__34001\,
            in3 => \N__34769\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => 'H',
            sr => \N__47360\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34768\,
            in2 => \_gnd_net_\,
            in3 => \N__32361\,
            lcout => \phase_controller_inst2.time_passed_RNI9M3O\,
            ltout => \phase_controller_inst2.time_passed_RNI9M3O_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_3_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__32399\,
            in1 => \N__32084\,
            in2 => \N__32048\,
            in3 => \N__37585\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => 'H',
            sr => \N__47360\
        );

    \phase_controller_inst2.start_timer_tr_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__34812\,
            in1 => \N__32045\,
            in2 => \N__34677\,
            in3 => \N__33962\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => 'H',
            sr => \N__47367\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34660\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => 'H',
            sr => \N__47367\
        );

    \phase_controller_inst2.T23_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__32023\,
            in1 => \N__34036\,
            in2 => \_gnd_net_\,
            in3 => \N__32368\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47768\,
            ce => 'H',
            sr => \N__47376\
        );

    \phase_controller_inst2.T45_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__32408\,
            in1 => \N__32335\,
            in2 => \_gnd_net_\,
            in3 => \N__32369\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47768\,
            ce => 'H',
            sr => \N__47376\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36407\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34147\,
            in2 => \_gnd_net_\,
            in3 => \N__34802\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47763\,
            ce => 'H',
            sr => \N__47383\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__32218\,
            in1 => \N__32275\,
            in2 => \_gnd_net_\,
            in3 => \N__32244\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_433_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__32219\,
            in1 => \N__32276\,
            in2 => \_gnd_net_\,
            in3 => \N__32245\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47758\,
            ce => 'H',
            sr => \N__47405\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32600\,
            in1 => \N__34059\,
            in2 => \_gnd_net_\,
            in3 => \N__32195\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_5_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__47855\,
            ce => \N__33335\,
            sr => \N__47285\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32596\,
            in1 => \N__34338\,
            in2 => \_gnd_net_\,
            in3 => \N__32192\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__47855\,
            ce => \N__33335\,
            sr => \N__47285\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32601\,
            in1 => \N__32835\,
            in2 => \_gnd_net_\,
            in3 => \N__32189\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__47855\,
            ce => \N__33335\,
            sr => \N__47285\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32597\,
            in1 => \N__32809\,
            in2 => \_gnd_net_\,
            in3 => \N__32186\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__47855\,
            ce => \N__33335\,
            sr => \N__47285\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32602\,
            in1 => \N__32784\,
            in2 => \_gnd_net_\,
            in3 => \N__32447\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__47855\,
            ce => \N__33335\,
            sr => \N__47285\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32598\,
            in1 => \N__32760\,
            in2 => \_gnd_net_\,
            in3 => \N__32444\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__47855\,
            ce => \N__33335\,
            sr => \N__47285\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32603\,
            in1 => \N__32731\,
            in2 => \_gnd_net_\,
            in3 => \N__32441\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__47855\,
            ce => \N__33335\,
            sr => \N__47285\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32599\,
            in1 => \N__32701\,
            in2 => \_gnd_net_\,
            in3 => \N__32438\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__47855\,
            ce => \N__33335\,
            sr => \N__47285\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32591\,
            in1 => \N__32673\,
            in2 => \_gnd_net_\,
            in3 => \N__32435\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__47844\,
            ce => \N__33338\,
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32595\,
            in1 => \N__32643\,
            in2 => \_gnd_net_\,
            in3 => \N__32432\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__47844\,
            ce => \N__33338\,
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32588\,
            in1 => \N__33061\,
            in2 => \_gnd_net_\,
            in3 => \N__32429\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__47844\,
            ce => \N__33338\,
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32592\,
            in1 => \N__33037\,
            in2 => \_gnd_net_\,
            in3 => \N__32426\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__47844\,
            ce => \N__33338\,
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32589\,
            in1 => \N__33012\,
            in2 => \_gnd_net_\,
            in3 => \N__32423\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__47844\,
            ce => \N__33338\,
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32593\,
            in1 => \N__32985\,
            in2 => \_gnd_net_\,
            in3 => \N__32474\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__47844\,
            ce => \N__33338\,
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32590\,
            in1 => \N__32959\,
            in2 => \_gnd_net_\,
            in3 => \N__32471\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__47844\,
            ce => \N__33338\,
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32594\,
            in1 => \N__32931\,
            in2 => \_gnd_net_\,
            in3 => \N__32468\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__47844\,
            ce => \N__33338\,
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32560\,
            in1 => \N__32901\,
            in2 => \_gnd_net_\,
            in3 => \N__32465\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__47835\,
            ce => \N__33337\,
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32564\,
            in1 => \N__32871\,
            in2 => \_gnd_net_\,
            in3 => \N__32462\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__47835\,
            ce => \N__33337\,
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32561\,
            in1 => \N__33279\,
            in2 => \_gnd_net_\,
            in3 => \N__32459\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__47835\,
            ce => \N__33337\,
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32565\,
            in1 => \N__33258\,
            in2 => \_gnd_net_\,
            in3 => \N__32456\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__47835\,
            ce => \N__33337\,
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32562\,
            in1 => \N__33231\,
            in2 => \_gnd_net_\,
            in3 => \N__32453\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__47835\,
            ce => \N__33337\,
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32566\,
            in1 => \N__33204\,
            in2 => \_gnd_net_\,
            in3 => \N__32450\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__47835\,
            ce => \N__33337\,
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32563\,
            in1 => \N__33178\,
            in2 => \_gnd_net_\,
            in3 => \N__32624\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__47835\,
            ce => \N__33337\,
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32567\,
            in1 => \N__33150\,
            in2 => \_gnd_net_\,
            in3 => \N__32621\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__47835\,
            ce => \N__33337\,
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32556\,
            in1 => \N__33117\,
            in2 => \_gnd_net_\,
            in3 => \N__32618\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__47828\,
            ce => \N__33336\,
            sr => \N__47305\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32568\,
            in1 => \N__33093\,
            in2 => \_gnd_net_\,
            in3 => \N__32615\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__47828\,
            ce => \N__33336\,
            sr => \N__47305\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32557\,
            in1 => \N__33462\,
            in2 => \_gnd_net_\,
            in3 => \N__32612\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__47828\,
            ce => \N__33336\,
            sr => \N__47305\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32569\,
            in1 => \N__33399\,
            in2 => \_gnd_net_\,
            in3 => \N__32609\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__47828\,
            ce => \N__33336\,
            sr => \N__47305\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32558\,
            in1 => \N__33442\,
            in2 => \_gnd_net_\,
            in3 => \N__32606\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__47828\,
            ce => \N__33336\,
            sr => \N__47305\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__33424\,
            in1 => \N__32559\,
            in2 => \_gnd_net_\,
            in3 => \N__32477\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47828\,
            ce => \N__33336\,
            sr => \N__47305\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34064\,
            in2 => \N__32846\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47823\,
            ce => \N__34300\,
            sr => \N__47311\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32815\,
            in2 => \N__34352\,
            in3 => \N__32849\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47823\,
            ce => \N__34300\,
            sr => \N__47311\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32845\,
            in2 => \N__32791\,
            in3 => \N__32819\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47823\,
            ce => \N__34300\,
            sr => \N__47311\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32816\,
            in2 => \N__32765\,
            in3 => \N__32795\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47823\,
            ce => \N__34300\,
            sr => \N__47311\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32737\,
            in2 => \N__32792\,
            in3 => \N__32768\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47823\,
            ce => \N__34300\,
            sr => \N__47311\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32764\,
            in2 => \N__32713\,
            in3 => \N__32741\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47823\,
            ce => \N__34300\,
            sr => \N__47311\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32738\,
            in2 => \N__32680\,
            in3 => \N__32717\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47823\,
            ce => \N__34300\,
            sr => \N__47311\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32644\,
            in2 => \N__32714\,
            in3 => \N__32687\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47823\,
            ce => \N__34300\,
            sr => \N__47311\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33067\,
            in2 => \N__32684\,
            in3 => \N__32654\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47818\,
            ce => \N__34302\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33043\,
            in2 => \N__32651\,
            in3 => \N__33071\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47818\,
            ce => \N__34302\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33068\,
            in2 => \N__33019\,
            in3 => \N__33047\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47818\,
            ce => \N__34302\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33044\,
            in2 => \N__32992\,
            in3 => \N__33023\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47818\,
            ce => \N__34302\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32965\,
            in2 => \N__33020\,
            in3 => \N__32996\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47818\,
            ce => \N__34302\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32938\,
            in2 => \N__32993\,
            in3 => \N__32969\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47818\,
            ce => \N__34302\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32966\,
            in2 => \N__32908\,
            in3 => \N__32945\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47818\,
            ce => \N__34302\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32872\,
            in2 => \N__32942\,
            in3 => \N__32915\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47818\,
            ce => \N__34302\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33280\,
            in2 => \N__32912\,
            in3 => \N__32882\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47812\,
            ce => \N__34303\,
            sr => \N__47319\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33259\,
            in2 => \N__32879\,
            in3 => \N__32852\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47812\,
            ce => \N__34303\,
            sr => \N__47319\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33281\,
            in2 => \N__33238\,
            in3 => \N__33263\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47812\,
            ce => \N__34303\,
            sr => \N__47319\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33260\,
            in2 => \N__33211\,
            in3 => \N__33242\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47812\,
            ce => \N__34303\,
            sr => \N__47319\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33184\,
            in2 => \N__33239\,
            in3 => \N__33215\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47812\,
            ce => \N__34303\,
            sr => \N__47319\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33157\,
            in2 => \N__33212\,
            in3 => \N__33188\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47812\,
            ce => \N__34303\,
            sr => \N__47319\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33185\,
            in2 => \N__33130\,
            in3 => \N__33164\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47812\,
            ce => \N__34303\,
            sr => \N__47319\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33094\,
            in2 => \N__33161\,
            in3 => \N__33134\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47812\,
            ce => \N__34303\,
            sr => \N__47319\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33463\,
            in2 => \N__33131\,
            in3 => \N__33101\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47806\,
            ce => \N__34304\,
            sr => \N__47324\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33406\,
            in2 => \N__33098\,
            in3 => \N__33074\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47806\,
            ce => \N__34304\,
            sr => \N__47324\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33464\,
            in2 => \N__33446\,
            in3 => \N__33428\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47806\,
            ce => \N__34304\,
            sr => \N__47324\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33425\,
            in2 => \N__33410\,
            in3 => \N__33383\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47806\,
            ce => \N__34304\,
            sr => \N__47324\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33380\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47806\,
            ce => \N__34304\,
            sr => \N__47324\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__33366\,
            in1 => \N__33840\,
            in2 => \_gnd_net_\,
            in3 => \N__33815\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_435_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36437\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__34719\,
            in1 => \N__34734\,
            in2 => \_gnd_net_\,
            in3 => \N__34678\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQ1_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33287\,
            in3 => \N__34612\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNI2FGQZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__34720\,
            in1 => \N__34679\,
            in2 => \_gnd_net_\,
            in3 => \N__35546\,
            lcout => \phase_controller_inst2.stoper_tr.running_1_sqmuxa\,
            ltout => \phase_controller_inst2.stoper_tr.running_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__34735\,
            in1 => \N__34680\,
            in2 => \N__33284\,
            in3 => \N__34721\,
            lcout => \phase_controller_inst2.stoper_tr.un1_start_latched2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33820\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33797\,
            ce => 'H',
            sr => \N__47331\
        );

    \delay_measurement_inst.start_timer_tr_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33819\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33797\,
            ce => 'H',
            sr => \N__47331\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36467\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33691\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44586\,
            in1 => \N__48084\,
            in2 => \N__45070\,
            in3 => \N__41111\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44626\,
            in1 => \N__45237\,
            in2 => \N__45488\,
            in3 => \N__43882\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36422\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44628\,
            in1 => \N__45234\,
            in2 => \N__46361\,
            in3 => \N__43613\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__45233\,
            in1 => \N__44627\,
            in2 => \N__41216\,
            in3 => \N__46424\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44625\,
            in1 => \N__45236\,
            in2 => \N__45917\,
            in3 => \N__40774\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45235\,
            in1 => \N__44629\,
            in2 => \N__46241\,
            in3 => \N__43552\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__38798\,
            in1 => \N__38557\,
            in2 => \_gnd_net_\,
            in3 => \N__34091\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__40637\,
            in1 => \_gnd_net_\,
            in2 => \N__33866\,
            in3 => \N__38799\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__46873\,
            in1 => \N__44622\,
            in2 => \N__41002\,
            in3 => \N__45241\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44623\,
            in1 => \N__48242\,
            in2 => \N__45278\,
            in3 => \N__45323\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36664\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44025\,
            in1 => \N__46872\,
            in2 => \_gnd_net_\,
            in3 => \N__40995\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44014\,
            in1 => \N__46234\,
            in2 => \_gnd_net_\,
            in3 => \N__43553\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44621\,
            in1 => \N__45915\,
            in2 => \N__45279\,
            in3 => \N__40778\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44624\,
            in1 => \N__46874\,
            in2 => \N__45280\,
            in3 => \N__41003\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43996\,
            in1 => \N__46946\,
            in2 => \_gnd_net_\,
            in3 => \N__41156\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34026\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34000\,
            lcout => \phase_controller_inst2.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36497\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011011100"
        )
    port map (
            in0 => \N__36980\,
            in1 => \N__35930\,
            in2 => \N__33941\,
            in3 => \N__33902\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44657\,
            in1 => \N__48002\,
            in2 => \N__41288\,
            in3 => \N__45147\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_1_11_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__45146\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44658\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44655\,
            in1 => \N__46750\,
            in2 => \N__40970\,
            in3 => \N__45148\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__46751\,
            in1 => \N__40969\,
            in2 => \N__45232\,
            in3 => \N__44656\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43997\,
            in1 => \N__46749\,
            in2 => \_gnd_net_\,
            in3 => \N__40965\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47021\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47773\,
            ce => \N__47509\,
            sr => \N__47368\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44659\,
            in1 => \N__48167\,
            in2 => \N__45293\,
            in3 => \N__44201\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44660\,
            in1 => \N__48001\,
            in2 => \N__45292\,
            in3 => \N__41284\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34146\,
            in2 => \_gnd_net_\,
            in3 => \N__34801\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47020\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47760\,
            ce => \N__47508\,
            sr => \N__47400\
        );

    \phase_controller_inst1.S2_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38438\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47759\,
            ce => 'H',
            sr => \N__47406\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34063\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47856\,
            ce => \N__34299\,
            sr => \N__47286\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__34404\,
            in1 => \N__34474\,
            in2 => \N__34448\,
            in3 => \N__34181\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_359_1\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_359_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__47470\,
            in1 => \N__34230\,
            in2 => \N__34184\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34318\,
            in1 => \N__41896\,
            in2 => \N__34367\,
            in3 => \N__37392\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_345\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__35386\,
            in1 => \N__37720\,
            in2 => \N__34175\,
            in3 => \N__35200\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__39574\,
            in1 => \N__41820\,
            in2 => \N__40079\,
            in3 => \N__34319\,
            lcout => \elapsed_time_ns_1_RNIAE2591_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__34475\,
            in1 => \N__34446\,
            in2 => \N__34253\,
            in3 => \N__34405\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40127\,
            in1 => \N__34271\,
            in2 => \N__37903\,
            in3 => \N__35193\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34207\,
            in1 => \N__37687\,
            in2 => \N__35107\,
            in3 => \N__41877\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__35103\,
            in1 => \N__34208\,
            in2 => \N__37393\,
            in3 => \N__34317\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__34169\,
            in1 => \N__41878\,
            in2 => \N__34172\,
            in3 => \N__34366\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37686\,
            in1 => \N__40131\,
            in2 => \N__37902\,
            in3 => \N__35192\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35119\,
            in2 => \_gnd_net_\,
            in3 => \N__37657\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34351\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47836\,
            ce => \N__34301\,
            sr => \N__47301\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__40132\,
            in1 => \N__34457\,
            in2 => \_gnd_net_\,
            in3 => \N__34280\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_349_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__40096\,
            in1 => \N__34270\,
            in2 => \N__34259\,
            in3 => \N__37889\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__38167\,
            in1 => \N__34406\,
            in2 => \N__34256\,
            in3 => \N__34473\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__34447\,
            in1 => \N__34252\,
            in2 => \N__34238\,
            in3 => \N__47471\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__47472\,
            in1 => \N__34232\,
            in2 => \N__34235\,
            in3 => \N__38170\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__34231\,
            in1 => \N__34217\,
            in2 => \N__35153\,
            in3 => \N__38168\,
            lcout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\,
            ltout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__38245\,
            in1 => \N__34201\,
            in2 => \N__34187\,
            in3 => \N__41555\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__35222\,
            in1 => \N__34424\,
            in2 => \N__41754\,
            in3 => \N__40038\,
            lcout => \elapsed_time_ns_1_RNI1HIF91_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__40039\,
            in1 => \N__34484\,
            in2 => \N__41769\,
            in3 => \N__37963\,
            lcout => \elapsed_time_ns_1_RNIQ9IF91_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__41700\,
            in1 => \N__35447\,
            in2 => \N__40068\,
            in3 => \N__34498\,
            lcout => \elapsed_time_ns_1_RNI0GIF91_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35239\,
            in1 => \N__34373\,
            in2 => \N__34499\,
            in3 => \N__34483\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35356\,
            in1 => \N__35398\,
            in2 => \N__35335\,
            in3 => \N__35278\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_347\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__40095\,
            in1 => \N__35382\,
            in2 => \N__34451\,
            in3 => \N__37716\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__34535\,
            in1 => \N__34385\,
            in2 => \N__41753\,
            in3 => \N__40037\,
            lcout => \elapsed_time_ns_1_RNIUDIF91_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35257\,
            in1 => \N__35425\,
            in2 => \N__34423\,
            in3 => \N__35164\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38014\,
            in1 => \N__38032\,
            in2 => \N__34562\,
            in3 => \N__34384\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36452\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__41721\,
            in1 => \N__34561\,
            in2 => \N__34547\,
            in3 => \N__40052\,
            lcout => \elapsed_time_ns_1_RNITCIF91_0_23\,
            ltout => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34538\,
            in3 => \N__34534\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36482\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34509\,
            in2 => \_gnd_net_\,
            in3 => \N__36189\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__37484\,
            in1 => \N__34828\,
            in2 => \N__34514\,
            in3 => \N__36220\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47813\,
            ce => 'H',
            sr => \N__47320\
        );

    \phase_controller_inst1.state_2_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__37520\,
            in1 => \N__34510\,
            in2 => \N__37565\,
            in3 => \N__36190\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47813\,
            ce => 'H',
            sr => \N__47320\
        );

    \phase_controller_inst1.state_1_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__34511\,
            in1 => \N__36191\,
            in2 => \N__38427\,
            in3 => \N__38395\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47813\,
            ce => 'H',
            sr => \N__47320\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38417\,
            in2 => \_gnd_net_\,
            in3 => \N__38394\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__38353\,
            in1 => \N__43020\,
            in2 => \N__34832\,
            in3 => \N__34829\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47813\,
            ce => 'H',
            sr => \N__47320\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__42958\,
            in1 => \N__42907\,
            in2 => \_gnd_net_\,
            in3 => \N__43016\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__34682\,
            in1 => \N__34761\,
            in2 => \N__34778\,
            in3 => \N__34717\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47807\,
            ce => 'H',
            sr => \N__47325\
        );

    \phase_controller_inst2.stoper_tr.running_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001010101110"
        )
    port map (
            in0 => \N__34736\,
            in1 => \N__34585\,
            in2 => \N__34745\,
            in3 => \N__34718\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47807\,
            ce => 'H',
            sr => \N__47325\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIP8O21_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__34716\,
            in1 => \N__34681\,
            in2 => \_gnd_net_\,
            in3 => \N__35539\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34601\,
            in3 => \N__34584\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34963\,
            in2 => \N__38324\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43797\,
            in2 => \N__43835\,
            in3 => \N__38577\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38578\,
            in1 => \N__44848\,
            in2 => \N__40679\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34859\,
            in2 => \N__45041\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44852\,
            in2 => \N__38309\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38297\,
            in2 => \N__45042\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44856\,
            in2 => \N__38477\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38486\,
            in2 => \N__45043\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38447\,
            in2 => \N__45044\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44863\,
            in2 => \N__34850\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43895\,
            in2 => \N__45045\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44867\,
            in2 => \N__34841\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34877\,
            in2 => \N__45046\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44871\,
            in2 => \N__45401\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34871\,
            in2 => \N__45047\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44875\,
            in2 => \N__43475\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44964\,
            in2 => \N__43199\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43625\,
            in2 => \N__45132\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44968\,
            in2 => \N__41129\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34865\,
            in2 => \N__45133\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44972\,
            in2 => \N__36650\,
            in3 => \N__34940\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34937\,
            in2 => \N__45134\,
            in3 => \N__34928\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44976\,
            in2 => \N__36623\,
            in3 => \N__34925\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36614\,
            in2 => \N__45135\,
            in3 => \N__34922\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45010\,
            in2 => \N__45347\,
            in3 => \N__34919\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34916\,
            in2 => \N__45143\,
            in3 => \N__34910\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45014\,
            in2 => \N__44177\,
            in3 => \N__34907\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34904\,
            in2 => \N__45144\,
            in3 => \N__34895\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45018\,
            in2 => \N__34892\,
            in3 => \N__34880\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44129\,
            in2 => \N__45145\,
            in3 => \N__34982\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45022\,
            in2 => \N__44243\,
            in3 => \N__34979\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_0_11_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010100110101"
        )
    port map (
            in0 => \N__35027\,
            in1 => \N__34976\,
            in2 => \N__38747\,
            in3 => \N__34967\,
            lcout => \current_shift_inst.control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34964\,
            in2 => \N__40636\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43801\,
            in2 => \N__43778\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44936\,
            in2 => \N__40664\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34946\,
            in2 => \N__45125\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44940\,
            in2 => \N__43232\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38498\,
            in2 => \N__45126\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44944\,
            in2 => \N__38465\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38270\,
            in2 => \N__45127\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44948\,
            in2 => \N__38288\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41225\,
            in2 => \N__45128\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44952\,
            in2 => \N__44114\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37277\,
            in2 => \N__45129\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44956\,
            in2 => \N__43586\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41297\,
            in2 => \N__45130\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44960\,
            in2 => \N__43526\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37262\,
            in2 => \N__45131\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37283\,
            in2 => \N__45136\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44983\,
            in2 => \N__37271\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41039\,
            in2 => \N__45137\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44987\,
            in2 => \N__35018\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36767\,
            in2 => \N__45138\,
            in3 => \N__35003\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44991\,
            in2 => \N__35000\,
            in3 => \N__34991\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39098\,
            in2 => \N__45139\,
            in3 => \N__34988\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44995\,
            in2 => \N__37637\,
            in3 => \N__34985\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44996\,
            in2 => \N__45446\,
            in3 => \N__35069\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44306\,
            in2 => \N__45140\,
            in3 => \N__35066\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45000\,
            in2 => \N__35063\,
            in3 => \N__35054\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40409\,
            in2 => \N__45141\,
            in3 => \N__35051\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45004\,
            in2 => \N__35048\,
            in3 => \N__35039\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39110\,
            in2 => \N__45142\,
            in3 => \N__35036\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45008\,
            in2 => \N__44242\,
            in3 => \N__35033\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_2_11_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__45009\,
            in1 => \N__44646\,
            in2 => \_gnd_net_\,
            in3 => \N__35030\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S1_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37551\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47765\,
            ce => 'H',
            sr => \N__47384\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001110"
        )
    port map (
            in0 => \N__42695\,
            in1 => \N__41582\,
            in2 => \N__41821\,
            in3 => \N__35207\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__35174\,
            in1 => \N__37996\,
            in2 => \N__41825\,
            in3 => \N__40076\,
            lcout => \elapsed_time_ns_1_RNIRBJF91_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42154\,
            in2 => \_gnd_net_\,
            in3 => \N__39564\,
            lcout => \phase_controller_inst1.stoper_tr.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__47469\,
            in1 => \N__35146\,
            in2 => \N__38174\,
            in3 => \N__35135\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__41516\,
            in1 => \_gnd_net_\,
            in2 => \N__35129\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIFG4DM1_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__40077\,
            in1 => \N__42366\,
            in2 => \N__41796\,
            in3 => \N__35126\,
            lcout => \elapsed_time_ns_1_RNIDH2591_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35075\,
            in2 => \_gnd_net_\,
            in3 => \N__41496\,
            lcout => \elapsed_time_ns_1_RNIIJ4DM1_0_19\,
            ltout => \elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__41743\,
            in1 => \N__35108\,
            in2 => \N__35078\,
            in3 => \N__41561\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__38093\,
            in1 => \N__42527\,
            in2 => \N__39896\,
            in3 => \N__39735\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47845\,
            ce => \N__43373\,
            sr => \N__47294\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__42523\,
            in1 => \N__37769\,
            in2 => \N__39764\,
            in3 => \N__38094\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47845\,
            ce => \N__43373\,
            sr => \N__47294\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__38091\,
            in1 => \N__42525\,
            in2 => \N__37799\,
            in3 => \N__39742\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47845\,
            ce => \N__43373\,
            sr => \N__47294\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__35285\,
            in1 => \N__37816\,
            in2 => \N__41768\,
            in3 => \N__40045\,
            lcout => \elapsed_time_ns_1_RNISAHF91_0_13\,
            ltout => \elapsed_time_ns_1_RNISAHF91_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__38092\,
            in1 => \N__42526\,
            in2 => \N__35267\,
            in3 => \N__39734\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47845\,
            ce => \N__43373\,
            sr => \N__47294\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__42524\,
            in1 => \N__37743\,
            in2 => \N__39765\,
            in3 => \N__38095\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47845\,
            ce => \N__43373\,
            sr => \N__47294\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__39732\,
            in1 => \N__42528\,
            in2 => \_gnd_net_\,
            in3 => \N__39271\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47845\,
            ce => \N__43373\,
            sr => \N__47294\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__42529\,
            in1 => \N__38246\,
            in2 => \_gnd_net_\,
            in3 => \N__39733\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47845\,
            ce => \N__43373\,
            sr => \N__47294\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__40035\,
            in1 => \N__35264\,
            in2 => \N__41770\,
            in3 => \N__37982\,
            lcout => \elapsed_time_ns_1_RNI3JIF91_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__35246\,
            in1 => \N__35228\,
            in2 => \N__41750\,
            in3 => \N__40030\,
            lcout => \elapsed_time_ns_1_RNIVEIF91_0_25\,
            ltout => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35413\,
            in1 => \N__35221\,
            in2 => \N__35210\,
            in3 => \N__35446\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__41685\,
            in1 => \N__35414\,
            in2 => \N__35435\,
            in3 => \N__40032\,
            lcout => \elapsed_time_ns_1_RNI2IIF91_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__40031\,
            in1 => \N__41689\,
            in2 => \N__35405\,
            in3 => \N__37771\,
            lcout => \elapsed_time_ns_1_RNIP7HF91_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__39513\,
            in1 => \N__35387\,
            in2 => \N__41752\,
            in3 => \N__40036\,
            lcout => \elapsed_time_ns_1_RNIGK2591_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__40033\,
            in1 => \N__41690\,
            in2 => \N__35363\,
            in3 => \N__37745\,
            lcout => \elapsed_time_ns_1_RNIR9HF91_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__37798\,
            in1 => \N__35339\,
            in2 => \N__41751\,
            in3 => \N__40034\,
            lcout => \elapsed_time_ns_1_RNIQ8HF91_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39629\,
            in2 => \N__35318\,
            in3 => \N__35755\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39599\,
            in2 => \N__35309\,
            in3 => \N__35717\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42128\,
            in2 => \N__35297\,
            in3 => \N__35687\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35528\,
            in2 => \N__42551\,
            in3 => \N__35669\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42344\,
            in2 => \N__35522\,
            in3 => \N__35651\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35633\,
            in1 => \N__39455\,
            in2 => \N__35510\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39209\,
            in2 => \N__35498\,
            in3 => \N__36110\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39611\,
            in2 => \N__35489\,
            in3 => \N__36092\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38048\,
            in2 => \N__35477\,
            in3 => \N__36074\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37862\,
            in2 => \N__35468\,
            in3 => \N__36056\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36038\,
            in1 => \N__35459\,
            in2 => \N__37850\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35453\,
            in2 => \N__37838\,
            in3 => \N__36020\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37826\,
            in2 => \N__35615\,
            in3 => \N__36002\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35981\,
            in1 => \N__37916\,
            in2 => \N__35606\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39221\,
            in2 => \N__35594\,
            in3 => \N__35963\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39236\,
            in2 => \N__35585\,
            in3 => \N__36392\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36374\,
            in1 => \N__38180\,
            in2 => \N__35576\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38210\,
            in2 => \N__35567\,
            in3 => \N__36356\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39251\,
            in2 => \N__35558\,
            in3 => \N__36335\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35549\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111101010"
        )
    port map (
            in0 => \N__35929\,
            in1 => \N__36944\,
            in2 => \N__35855\,
            in3 => \N__35822\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35765\,
            in2 => \N__35759\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42069\,
            in1 => \N__35716\,
            in2 => \_gnd_net_\,
            in3 => \N__35702\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__47814\,
            ce => 'H',
            sr => \N__47321\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__42081\,
            in1 => \N__35686\,
            in2 => \N__35699\,
            in3 => \N__35672\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__47814\,
            ce => 'H',
            sr => \N__47321\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42070\,
            in1 => \N__35668\,
            in2 => \_gnd_net_\,
            in3 => \N__35654\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__47814\,
            ce => 'H',
            sr => \N__47321\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42082\,
            in1 => \N__35650\,
            in2 => \_gnd_net_\,
            in3 => \N__35636\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__47814\,
            ce => 'H',
            sr => \N__47321\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42071\,
            in1 => \N__35632\,
            in2 => \_gnd_net_\,
            in3 => \N__35618\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__47814\,
            ce => 'H',
            sr => \N__47321\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42083\,
            in1 => \N__36109\,
            in2 => \_gnd_net_\,
            in3 => \N__36095\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__47814\,
            ce => 'H',
            sr => \N__47321\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42072\,
            in1 => \N__36091\,
            in2 => \_gnd_net_\,
            in3 => \N__36077\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__47814\,
            ce => 'H',
            sr => \N__47321\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42097\,
            in1 => \N__36073\,
            in2 => \_gnd_net_\,
            in3 => \N__36059\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__47808\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42089\,
            in1 => \N__36055\,
            in2 => \_gnd_net_\,
            in3 => \N__36041\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__47808\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42094\,
            in1 => \N__36037\,
            in2 => \_gnd_net_\,
            in3 => \N__36023\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__47808\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42090\,
            in1 => \N__36019\,
            in2 => \_gnd_net_\,
            in3 => \N__36005\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__47808\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42095\,
            in1 => \N__35998\,
            in2 => \_gnd_net_\,
            in3 => \N__35984\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__47808\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42091\,
            in1 => \N__35980\,
            in2 => \_gnd_net_\,
            in3 => \N__35966\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__47808\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42096\,
            in1 => \N__35959\,
            in2 => \_gnd_net_\,
            in3 => \N__35945\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__47808\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42092\,
            in1 => \N__36391\,
            in2 => \_gnd_net_\,
            in3 => \N__36377\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__47808\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42087\,
            in1 => \N__36373\,
            in2 => \_gnd_net_\,
            in3 => \N__36359\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__47802\,
            ce => 'H',
            sr => \N__47329\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42093\,
            in1 => \N__36355\,
            in2 => \_gnd_net_\,
            in3 => \N__36341\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__47802\,
            ce => 'H',
            sr => \N__47329\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42088\,
            in1 => \N__36334\,
            in2 => \_gnd_net_\,
            in3 => \N__36338\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47802\,
            ce => 'H',
            sr => \N__47329\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__36320\,
            in1 => \N__36308\,
            in2 => \N__36251\,
            in3 => \N__36180\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47802\,
            ce => 'H',
            sr => \N__47329\
        );

    \current_shift_inst.control_input_0_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36779\,
            in2 => \N__36638\,
            in3 => \N__36637\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__47796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36746\,
            in3 => \N__36128\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__47796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36719\,
            in2 => \_gnd_net_\,
            in3 => \N__36113\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__47796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36692\,
            in2 => \_gnd_net_\,
            in3 => \N__36500\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__47796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37349\,
            in2 => \_gnd_net_\,
            in3 => \N__36485\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__47796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37322\,
            in2 => \_gnd_net_\,
            in3 => \N__36470\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__47796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37292\,
            in2 => \_gnd_net_\,
            in3 => \N__36455\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__47796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36593\,
            in2 => \_gnd_net_\,
            in3 => \N__36440\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__47796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36566\,
            in2 => \_gnd_net_\,
            in3 => \N__36425\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__47791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36542\,
            in2 => \_gnd_net_\,
            in3 => \N__36410\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__47791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36518\,
            in2 => \_gnd_net_\,
            in3 => \N__36395\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__47791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36683\,
            in2 => \_gnd_net_\,
            in3 => \N__36674\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44618\,
            in1 => \N__46817\,
            in2 => \N__45202\,
            in3 => \N__41071\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38740\,
            lcout => \current_shift_inst.N_1609_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44619\,
            in1 => \N__46692\,
            in2 => \N__45201\,
            in3 => \N__40942\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45098\,
            in1 => \N__44620\,
            in2 => \N__46628\,
            in3 => \N__40911\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__36608\,
            in1 => \N__36602\,
            in2 => \_gnd_net_\,
            in3 => \N__38733\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38734\,
            in1 => \N__36584\,
            in2 => \_gnd_net_\,
            in3 => \N__36572\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__36560\,
            in1 => \N__36554\,
            in2 => \_gnd_net_\,
            in3 => \N__38735\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38736\,
            in1 => \N__36536\,
            in2 => \_gnd_net_\,
            in3 => \N__36524\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__37157\,
            in1 => \N__36998\,
            in2 => \N__37200\,
            in3 => \N__37243\,
            lcout => \elapsed_time_ns_1_RNI81DJ11_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37229\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47786\,
            ce => \N__37178\,
            sr => \N__47339\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__37156\,
            in1 => \N__36808\,
            in2 => \N__37025\,
            in3 => \N__36997\,
            lcout => \elapsed_time_ns_1_RNIO1ND11_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__36794\,
            in1 => \N__36785\,
            in2 => \_gnd_net_\,
            in3 => \N__38723\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46813\,
            in1 => \N__44653\,
            in2 => \N__45263\,
            in3 => \N__41075\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__36761\,
            in1 => \N__38724\,
            in2 => \_gnd_net_\,
            in3 => \N__36752\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__38725\,
            in1 => \N__36734\,
            in2 => \_gnd_net_\,
            in3 => \N__36725\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__36707\,
            in1 => \N__36701\,
            in2 => \_gnd_net_\,
            in3 => \N__38726\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38728\,
            in1 => \N__37367\,
            in2 => \_gnd_net_\,
            in3 => \N__37358\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__37340\,
            in1 => \N__37331\,
            in2 => \_gnd_net_\,
            in3 => \N__38727\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__38729\,
            in1 => \_gnd_net_\,
            in2 => \N__37313\,
            in3 => \N__37301\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44649\,
            in1 => \N__45209\,
            in2 => \N__46112\,
            in3 => \N__43709\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44065\,
            in1 => \N__46693\,
            in2 => \_gnd_net_\,
            in3 => \N__40943\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__45207\,
            in1 => \N__44647\,
            in2 => \N__41215\,
            in3 => \N__46423\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44650\,
            in1 => \N__46054\,
            in2 => \N__43667\,
            in3 => \N__45210\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__46620\,
            in1 => \N__40912\,
            in2 => \_gnd_net_\,
            in3 => \N__44066\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44648\,
            in1 => \N__45208\,
            in2 => \N__46169\,
            in3 => \N__43504\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45206\,
            in1 => \N__44651\,
            in2 => \N__46627\,
            in3 => \N__40913\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__37543\,
            in1 => \N__37423\,
            in2 => \N__37459\,
            in3 => \N__37600\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47774\,
            ce => 'H',
            sr => \N__47369\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39142\,
            in2 => \_gnd_net_\,
            in3 => \N__37418\,
            lcout => \current_shift_inst.timer_s1.N_166_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.start_timer_s1_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__37599\,
            in1 => \N__37452\,
            in2 => \_gnd_net_\,
            in3 => \N__37547\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47774\,
            ce => 'H',
            sr => \N__47369\
        );

    \phase_controller_inst1.state_3_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__38357\,
            in1 => \N__37519\,
            in2 => \N__37552\,
            in3 => \N__37586\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47774\,
            ce => 'H',
            sr => \N__47369\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37542\,
            in2 => \_gnd_net_\,
            in3 => \N__37518\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__39143\,
            in1 => \N__37419\,
            in2 => \_gnd_net_\,
            in3 => \N__37451\,
            lcout => \current_shift_inst.timer_s1.N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__37469\,
            in1 => \N__39126\,
            in2 => \_gnd_net_\,
            in3 => \N__37433\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47866\,
            ce => 'H',
            sr => \N__47281\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__42164\,
            in1 => \N__41803\,
            in2 => \N__41497\,
            in3 => \N__37397\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__41584\,
            in1 => \_gnd_net_\,
            in2 => \N__37697\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIRHL2M1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101110"
        )
    port map (
            in0 => \N__38195\,
            in1 => \N__41583\,
            in2 => \N__37694\,
            in3 => \N__41804\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37670\,
            in3 => \N__41480\,
            lcout => \elapsed_time_ns_1_RNIGH4DM1_0_17\,
            ltout => \elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__38238\,
            in1 => \N__41845\,
            in2 => \N__37667\,
            in3 => \N__39269\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__42567\,
            in1 => \N__37664\,
            in2 => \N__41822\,
            in3 => \N__40075\,
            lcout => \elapsed_time_ns_1_RNICG2591_0_4\,
            ltout => \elapsed_time_ns_1_RNICG2591_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38196\,
            in1 => \N__41846\,
            in2 => \N__37646\,
            in3 => \N__42360\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__39270\,
            in1 => \N__38237\,
            in2 => \N__37643\,
            in3 => \N__39946\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37868\,
            in2 => \_gnd_net_\,
            in3 => \N__41479\,
            lcout => \elapsed_time_ns_1_RNIDE4DM1_0_14\,
            ltout => \elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39839\,
            in2 => \N__37640\,
            in3 => \N__39806\,
            lcout => \phase_controller_inst1.stoper_tr.N_241\,
            ltout => \phase_controller_inst1.stoper_tr.N_241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__42520\,
            in1 => \N__39892\,
            in2 => \N__37919\,
            in3 => \N__39754\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47857\,
            ce => \N__42116\,
            sr => \N__47287\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__41586\,
            in1 => \N__39891\,
            in2 => \N__37907\,
            in3 => \N__41809\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__42518\,
            in1 => \N__37770\,
            in2 => \N__38108\,
            in3 => \N__39752\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47857\,
            ce => \N__42116\,
            sr => \N__47287\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__38089\,
            in1 => \N__42521\,
            in2 => \N__39766\,
            in3 => \N__37797\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47857\,
            ce => \N__42116\,
            sr => \N__47287\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__42519\,
            in1 => \N__37744\,
            in2 => \N__38109\,
            in3 => \N__39753\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47857\,
            ce => \N__42116\,
            sr => \N__47287\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__38090\,
            in1 => \N__42522\,
            in2 => \N__39767\,
            in3 => \N__37817\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47857\,
            ce => \N__42116\,
            sr => \N__47287\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__39477\,
            in1 => \N__42452\,
            in2 => \N__39756\,
            in3 => \N__39551\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37815\,
            in1 => \N__37793\,
            in2 => \N__37772\,
            in3 => \N__37742\,
            lcout => \phase_controller_inst1.stoper_tr.N_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__37721\,
            in1 => \N__42621\,
            in2 => \N__41816\,
            in3 => \N__40059\,
            lcout => \elapsed_time_ns_1_RNIFJ2591_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__40058\,
            in1 => \N__37949\,
            in2 => \N__38042\,
            in3 => \N__41786\,
            lcout => \elapsed_time_ns_1_RNISBIF91_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__38021\,
            in1 => \N__38003\,
            in2 => \N__41815\,
            in3 => \N__40057\,
            lcout => \elapsed_time_ns_1_RNIRAIF91_0_21\,
            ltout => \elapsed_time_ns_1_RNIRAIF91_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37997\,
            in1 => \N__37981\,
            in2 => \N__37970\,
            in3 => \N__37967\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37948\,
            in1 => \N__37940\,
            in2 => \N__37934\,
            in3 => \N__37931\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__39755\,
            in1 => \N__38117\,
            in2 => \N__39925\,
            in3 => \N__38111\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47837\,
            ce => \N__43367\,
            sr => \N__47302\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__39743\,
            in1 => \N__42510\,
            in2 => \_gnd_net_\,
            in3 => \N__38204\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47837\,
            ce => \N__43367\,
            sr => \N__47302\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__41860\,
            in1 => \N__42450\,
            in2 => \_gnd_net_\,
            in3 => \N__39745\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47837\,
            ce => \N__43367\,
            sr => \N__47302\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__39744\,
            in1 => \N__39845\,
            in2 => \N__39811\,
            in3 => \N__42511\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47837\,
            ce => \N__43367\,
            sr => \N__47302\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__42289\,
            in1 => \N__42451\,
            in2 => \_gnd_net_\,
            in3 => \N__39509\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47837\,
            ce => \N__43367\,
            sr => \N__47302\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__42231\,
            in1 => \N__42290\,
            in2 => \N__42332\,
            in3 => \N__42169\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47837\,
            ce => \N__43367\,
            sr => \N__47302\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__39918\,
            in1 => \N__39802\,
            in2 => \_gnd_net_\,
            in3 => \N__39863\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38258\,
            in2 => \_gnd_net_\,
            in3 => \N__41504\,
            lcout => \elapsed_time_ns_1_RNIHI4DM1_0_18\,
            ltout => \elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__39758\,
            in1 => \_gnd_net_\,
            in2 => \N__38213\,
            in3 => \N__42433\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47829\,
            ce => \N__42119\,
            sr => \N__47306\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__42432\,
            in1 => \N__38203\,
            in2 => \_gnd_net_\,
            in3 => \N__39760\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47829\,
            ce => \N__42119\,
            sr => \N__47306\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__38169\,
            in1 => \N__42431\,
            in2 => \N__41823\,
            in3 => \N__40078\,
            lcout => \elapsed_time_ns_1_RNISCJF91_0_31\,
            ltout => \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111110"
        )
    port map (
            in0 => \N__38126\,
            in1 => \N__39950\,
            in2 => \N__38120\,
            in3 => \N__39757\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__39759\,
            in1 => \N__38110\,
            in2 => \N__38051\,
            in3 => \N__39926\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47829\,
            ce => \N__42119\,
            sr => \N__47306\
        );

    \phase_controller_inst1.state_0_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__38335\,
            in1 => \N__38428\,
            in2 => \N__38369\,
            in3 => \N__38399\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => 'H',
            sr => \N__47312\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38334\,
            in2 => \_gnd_net_\,
            in3 => \N__38365\,
            lcout => \phase_controller_inst1.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__38336\,
            in1 => \N__43024\,
            in2 => \N__42975\,
            in3 => \N__42878\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => 'H',
            sr => \N__47312\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43023\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => 'H',
            sr => \N__47312\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__42840\,
            in1 => \N__42865\,
            in2 => \N__42795\,
            in3 => \N__43351\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => 'H',
            sr => \N__47312\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__44417\,
            in1 => \N__40646\,
            in2 => \_gnd_net_\,
            in3 => \N__40480\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44426\,
            in1 => \N__45842\,
            in2 => \N__45176\,
            in3 => \N__43249\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44422\,
            in1 => \N__45051\,
            in2 => \N__45767\,
            in3 => \N__40732\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45061\,
            in1 => \N__44424\,
            in2 => \N__45548\,
            in3 => \N__40879\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44421\,
            in1 => \N__45060\,
            in2 => \N__45622\,
            in3 => \N__40697\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__40733\,
            in1 => \N__45763\,
            in2 => \N__45177\,
            in3 => \N__44420\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44423\,
            in1 => \N__45059\,
            in2 => \N__45623\,
            in3 => \N__40696\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44427\,
            in1 => \N__45691\,
            in2 => \N__45178\,
            in3 => \N__40714\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__40715\,
            in1 => \N__45058\,
            in2 => \N__45692\,
            in3 => \N__44425\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44081\,
            in1 => \N__45838\,
            in2 => \_gnd_net_\,
            in3 => \N__43248\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45916\,
            in1 => \N__44080\,
            in2 => \_gnd_net_\,
            in3 => \N__40762\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44534\,
            in1 => \N__45181\,
            in2 => \N__40880\,
            in3 => \N__45544\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45984\,
            in1 => \N__44079\,
            in2 => \_gnd_net_\,
            in3 => \N__40792\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44083\,
            in1 => \N__45682\,
            in2 => \_gnd_net_\,
            in3 => \N__40713\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45610\,
            in1 => \N__44084\,
            in2 => \_gnd_net_\,
            in3 => \N__40695\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44082\,
            in1 => \N__45757\,
            in2 => \_gnd_net_\,
            in3 => \N__40731\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45543\,
            in1 => \N__44085\,
            in2 => \_gnd_net_\,
            in3 => \N__40875\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38582\,
            in2 => \N__38558\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39035\,
            in2 => \N__43733\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38531\,
            in2 => \N__39064\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39039\,
            in2 => \N__38525\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38513\,
            in2 => \N__39065\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39043\,
            in2 => \N__38507\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38624\,
            in2 => \N__39066\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39047\,
            in2 => \N__38618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39030\,
            in2 => \N__38609\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39034\,
            in2 => \N__43856\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39027\,
            in2 => \N__43907\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39031\,
            in2 => \N__41177\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39028\,
            in2 => \N__41246\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39032\,
            in2 => \N__43568\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39029\,
            in2 => \N__38597\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39033\,
            in2 => \N__43214\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39011\,
            in2 => \N__43682\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41027\,
            in2 => \N__39060\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39015\,
            in2 => \N__38684\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38672\,
            in2 => \N__39061\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39019\,
            in2 => \N__41048\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38657\,
            in2 => \N__39062\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39023\,
            in2 => \N__38645\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38633\,
            in2 => \N__39063\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38850\,
            in2 => \N__41234\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44213\,
            in2 => \N__38922\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38854\,
            in2 => \N__41021\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40397\,
            in2 => \N__38923\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38858\,
            in2 => \N__41261\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41252\,
            in2 => \N__38924\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38862\,
            in2 => \N__44270\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44611\,
            in2 => \_gnd_net_\,
            in3 => \N__38750\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39141\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44654\,
            in1 => \N__47915\,
            in2 => \N__44159\,
            in3 => \N__45257\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44652\,
            in1 => \N__46694\,
            in2 => \N__45287\,
            in3 => \N__40941\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39402\,
            in1 => \N__46008\,
            in2 => \_gnd_net_\,
            in3 => \N__39089\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__47778\,
            ce => \N__39310\,
            sr => \N__47361\
        );

    \current_shift_inst.timer_s1.counter_1_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39406\,
            in1 => \N__45936\,
            in2 => \_gnd_net_\,
            in3 => \N__39086\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__47778\,
            ce => \N__39310\,
            sr => \N__47361\
        );

    \current_shift_inst.timer_s1.counter_2_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39403\,
            in1 => \N__45861\,
            in2 => \_gnd_net_\,
            in3 => \N__39083\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__47778\,
            ce => \N__39310\,
            sr => \N__47361\
        );

    \current_shift_inst.timer_s1.counter_3_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39407\,
            in1 => \N__45781\,
            in2 => \_gnd_net_\,
            in3 => \N__39080\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__47778\,
            ce => \N__39310\,
            sr => \N__47361\
        );

    \current_shift_inst.timer_s1.counter_4_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39404\,
            in1 => \N__45708\,
            in2 => \_gnd_net_\,
            in3 => \N__39077\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__47778\,
            ce => \N__39310\,
            sr => \N__47361\
        );

    \current_shift_inst.timer_s1.counter_5_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39408\,
            in1 => \N__45639\,
            in2 => \_gnd_net_\,
            in3 => \N__39074\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__47778\,
            ce => \N__39310\,
            sr => \N__47361\
        );

    \current_shift_inst.timer_s1.counter_6_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39405\,
            in1 => \N__45564\,
            in2 => \_gnd_net_\,
            in3 => \N__39071\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__47778\,
            ce => \N__39310\,
            sr => \N__47361\
        );

    \current_shift_inst.timer_s1.counter_7_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39409\,
            in1 => \N__45504\,
            in2 => \_gnd_net_\,
            in3 => \N__39170\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__47778\,
            ce => \N__39310\,
            sr => \N__47361\
        );

    \current_shift_inst.timer_s1.counter_8_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39421\,
            in1 => \N__46512\,
            in2 => \_gnd_net_\,
            in3 => \N__39167\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__47775\,
            ce => \N__39302\,
            sr => \N__47370\
        );

    \current_shift_inst.timer_s1.counter_9_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39431\,
            in1 => \N__46446\,
            in2 => \_gnd_net_\,
            in3 => \N__39164\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__47775\,
            ce => \N__39302\,
            sr => \N__47370\
        );

    \current_shift_inst.timer_s1.counter_10_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39418\,
            in1 => \N__46383\,
            in2 => \_gnd_net_\,
            in3 => \N__39161\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__47775\,
            ce => \N__39302\,
            sr => \N__47370\
        );

    \current_shift_inst.timer_s1.counter_11_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39428\,
            in1 => \N__46312\,
            in2 => \_gnd_net_\,
            in3 => \N__39158\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__47775\,
            ce => \N__39302\,
            sr => \N__47370\
        );

    \current_shift_inst.timer_s1.counter_12_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39419\,
            in1 => \N__46257\,
            in2 => \_gnd_net_\,
            in3 => \N__39155\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__47775\,
            ce => \N__39302\,
            sr => \N__47370\
        );

    \current_shift_inst.timer_s1.counter_13_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39429\,
            in1 => \N__46183\,
            in2 => \_gnd_net_\,
            in3 => \N__39152\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__47775\,
            ce => \N__39302\,
            sr => \N__47370\
        );

    \current_shift_inst.timer_s1.counter_14_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39420\,
            in1 => \N__46126\,
            in2 => \_gnd_net_\,
            in3 => \N__39149\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__47775\,
            ce => \N__39302\,
            sr => \N__47370\
        );

    \current_shift_inst.timer_s1.counter_15_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39430\,
            in1 => \N__46069\,
            in2 => \_gnd_net_\,
            in3 => \N__39146\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__47775\,
            ce => \N__39302\,
            sr => \N__47370\
        );

    \current_shift_inst.timer_s1.counter_16_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39410\,
            in1 => \N__46968\,
            in2 => \_gnd_net_\,
            in3 => \N__39197\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__47770\,
            ce => \N__39311\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.counter_17_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39422\,
            in1 => \N__46896\,
            in2 => \_gnd_net_\,
            in3 => \N__39194\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__47770\,
            ce => \N__39311\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.counter_18_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39411\,
            in1 => \N__46839\,
            in2 => \_gnd_net_\,
            in3 => \N__39191\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__47770\,
            ce => \N__39311\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.counter_19_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39423\,
            in1 => \N__46765\,
            in2 => \_gnd_net_\,
            in3 => \N__39188\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__47770\,
            ce => \N__39311\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.counter_20_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39412\,
            in1 => \N__46710\,
            in2 => \_gnd_net_\,
            in3 => \N__39185\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__47770\,
            ce => \N__39311\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.counter_21_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39424\,
            in1 => \N__46642\,
            in2 => \_gnd_net_\,
            in3 => \N__39182\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__47770\,
            ce => \N__39311\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.counter_22_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39413\,
            in1 => \N__46579\,
            in2 => \_gnd_net_\,
            in3 => \N__39179\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__47770\,
            ce => \N__39311\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.counter_23_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39425\,
            in1 => \N__48256\,
            in2 => \_gnd_net_\,
            in3 => \N__39176\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__47770\,
            ce => \N__39311\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.counter_24_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39414\,
            in1 => \N__48189\,
            in2 => \_gnd_net_\,
            in3 => \N__39173\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__47766\,
            ce => \N__39303\,
            sr => \N__47385\
        );

    \current_shift_inst.timer_s1.counter_25_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39426\,
            in1 => \N__48108\,
            in2 => \_gnd_net_\,
            in3 => \N__39443\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__47766\,
            ce => \N__39303\,
            sr => \N__47385\
        );

    \current_shift_inst.timer_s1.counter_26_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39415\,
            in1 => \N__48024\,
            in2 => \_gnd_net_\,
            in3 => \N__39440\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__47766\,
            ce => \N__39303\,
            sr => \N__47385\
        );

    \current_shift_inst.timer_s1.counter_27_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39427\,
            in1 => \N__47931\,
            in2 => \_gnd_net_\,
            in3 => \N__39437\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__47766\,
            ce => \N__39303\,
            sr => \N__47385\
        );

    \current_shift_inst.timer_s1.counter_28_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39416\,
            in1 => \N__48043\,
            in2 => \_gnd_net_\,
            in3 => \N__39434\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__47766\,
            ce => \N__39303\,
            sr => \N__47385\
        );

    \current_shift_inst.timer_s1.counter_29_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__47956\,
            in1 => \N__39417\,
            in2 => \_gnd_net_\,
            in3 => \N__39314\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47766\,
            ce => \N__39303\,
            sr => \N__47385\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__39761\,
            in1 => \N__42512\,
            in2 => \_gnd_net_\,
            in3 => \N__39275\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47867\,
            ce => \N__42117\,
            sr => \N__47282\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__42515\,
            in1 => \N__41856\,
            in2 => \_gnd_net_\,
            in3 => \N__39763\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47867\,
            ce => \N__42117\,
            sr => \N__47282\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__39762\,
            in1 => \N__39840\,
            in2 => \N__39815\,
            in3 => \N__42514\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47867\,
            ce => \N__42117\,
            sr => \N__47282\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__42516\,
            in1 => \N__42306\,
            in2 => \N__42626\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47867\,
            ce => \N__42117\,
            sr => \N__47282\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__42304\,
            in1 => \N__42513\,
            in2 => \_gnd_net_\,
            in3 => \N__39521\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47867\,
            ce => \N__42117\,
            sr => \N__47282\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__42517\,
            in1 => \N__42305\,
            in2 => \N__42239\,
            in3 => \N__42662\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47867\,
            ce => \N__42117\,
            sr => \N__47282\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__39714\,
            in1 => \N__39587\,
            in2 => \N__39482\,
            in3 => \N__39550\,
            lcout => \phase_controller_inst1.stoper_tr.N_235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101010101"
        )
    port map (
            in0 => \N__39575\,
            in1 => \N__39478\,
            in2 => \N__42165\,
            in3 => \N__39549\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41498\,
            in2 => \_gnd_net_\,
            in3 => \N__39533\,
            lcout => \elapsed_time_ns_1_RNIUKL2M1_0_6\,
            ltout => \elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__39520\,
            in1 => \N__42614\,
            in2 => \N__39485\,
            in3 => \N__39862\,
            lcout => \phase_controller_inst1.stoper_tr.N_247\,
            ltout => \phase_controller_inst1.stoper_tr.N_247_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39807\,
            in2 => \N__39461\,
            in3 => \N__39713\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__42690\,
            in1 => \N__42467\,
            in2 => \N__39458\,
            in3 => \N__42303\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47863\,
            ce => \N__42098\,
            sr => \N__47283\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101010"
        )
    port map (
            in0 => \N__41585\,
            in1 => \N__40133\,
            in2 => \N__41811\,
            in3 => \N__39917\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__40103\,
            in1 => \N__39800\,
            in2 => \N__41810\,
            in3 => \N__40056\,
            lcout => \elapsed_time_ns_1_RNIUCHF91_0_15\,
            ltout => \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39889\,
            in2 => \N__39953\,
            in3 => \N__39916\,
            lcout => \phase_controller_inst1.stoper_tr.N_251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39932\,
            in2 => \_gnd_net_\,
            in3 => \N__41499\,
            lcout => \elapsed_time_ns_1_RNI1OL2M1_0_9\,
            ltout => \elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39890\,
            in2 => \N__39866\,
            in3 => \N__39861\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.N_211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__39844\,
            in1 => \N__39801\,
            in2 => \N__39770\,
            in3 => \N__39715\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41430\,
            in2 => \N__39635\,
            in3 => \N__42453\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__41431\,
            in1 => \N__42224\,
            in2 => \N__39632\,
            in3 => \N__41413\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47858\,
            ce => \N__42118\,
            sr => \N__47288\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39617\,
            in2 => \N__41393\,
            in3 => \N__42796\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42647\,
            in2 => \N__40229\,
            in3 => \N__42763\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40220\,
            in2 => \N__40214\,
            in3 => \N__42739\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42641\,
            in2 => \N__40205\,
            in3 => \N__42724\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40196\,
            in2 => \N__42635\,
            in3 => \N__42709\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40190\,
            in2 => \N__42671\,
            in3 => \N__43180\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42593\,
            in2 => \N__40181\,
            in3 => \N__43165\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43150\,
            in1 => \N__40172\,
            in2 => \N__40160\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43135\,
            in1 => \N__40148\,
            in2 => \N__40142\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40370\,
            in2 => \N__40385\,
            in3 => \N__43120\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40364\,
            in2 => \N__40352\,
            in3 => \N__43105\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40343\,
            in2 => \N__40331\,
            in3 => \N__43090\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43075\,
            in1 => \N__40322\,
            in2 => \N__40310\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40286\,
            in2 => \N__40301\,
            in3 => \N__43447\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40280\,
            in2 => \N__40274\,
            in3 => \N__43432\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40265\,
            in2 => \N__40259\,
            in3 => \N__43417\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40250\,
            in2 => \N__40238\,
            in3 => \N__43402\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40454\,
            in2 => \N__40442\,
            in3 => \N__43387\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40433\,
            in2 => \N__40421\,
            in3 => \N__43261\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40412\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8I2_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42839\,
            in2 => \_gnd_net_\,
            in3 => \N__42864\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNISF8IZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__43022\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42945\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__43021\,
            in1 => \N__42944\,
            in2 => \_gnd_net_\,
            in3 => \N__43054\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000101"
        )
    port map (
            in0 => \N__48086\,
            in1 => \N__41107\,
            in2 => \N__44480\,
            in3 => \N__45198\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__41106\,
            in1 => \N__48085\,
            in2 => \_gnd_net_\,
            in3 => \N__44413\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47825\,
            ce => \N__47516\,
            sr => \N__47313\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45199\,
            in1 => \N__44412\,
            in2 => \N__45989\,
            in3 => \N__40798\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100011"
        )
    port map (
            in0 => \N__40799\,
            in1 => \N__45985\,
            in2 => \N__44479\,
            in3 => \N__45200\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40827\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44408\,
            in2 => \N__40640\,
            in3 => \N__40479\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40612\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40547\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40475\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46019\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47819\,
            ce => \N__47515\,
            sr => \N__47316\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45836\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45756\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43817\,
            in2 => \N__40828\,
            in3 => \N__40826\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43841\,
            in2 => \_gnd_net_\,
            in3 => \N__40781\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43460\,
            in2 => \_gnd_net_\,
            in3 => \N__40751\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40748\,
            in2 => \_gnd_net_\,
            in3 => \N__40742\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40739\,
            in2 => \_gnd_net_\,
            in3 => \N__40718\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44294\,
            in2 => \_gnd_net_\,
            in3 => \N__40700\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43454\,
            in2 => \_gnd_net_\,
            in3 => \N__40682\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44282\,
            in2 => \_gnd_net_\,
            in3 => \N__40862\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45383\,
            in2 => \_gnd_net_\,
            in3 => \N__40859\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41366\,
            in2 => \_gnd_net_\,
            in3 => \N__40856\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44165\,
            in2 => \_gnd_net_\,
            in3 => \N__40853\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41165\,
            in2 => \_gnd_net_\,
            in3 => \N__40850\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44120\,
            in2 => \_gnd_net_\,
            in3 => \N__40847\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41357\,
            in2 => \_gnd_net_\,
            in3 => \N__40844\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41324\,
            in2 => \_gnd_net_\,
            in3 => \N__40841\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41306\,
            in2 => \_gnd_net_\,
            in3 => \N__40838\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45374\,
            in2 => \_gnd_net_\,
            in3 => \N__41009\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41345\,
            in2 => \_gnd_net_\,
            in3 => \N__41006\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41384\,
            in2 => \_gnd_net_\,
            in3 => \N__40976\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43718\,
            in2 => \_gnd_net_\,
            in3 => \N__40973\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41375\,
            in2 => \_gnd_net_\,
            in3 => \N__40946\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45329\,
            in2 => \_gnd_net_\,
            in3 => \N__40916\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41942\,
            in2 => \_gnd_net_\,
            in3 => \N__40889\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41315\,
            in2 => \_gnd_net_\,
            in3 => \N__40886\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41951\,
            in2 => \_gnd_net_\,
            in3 => \N__40883\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41333\,
            in2 => \_gnd_net_\,
            in3 => \N__41114\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41915\,
            in2 => \_gnd_net_\,
            in3 => \N__41087\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41933\,
            in2 => \_gnd_net_\,
            in3 => \N__41084\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41924\,
            in2 => \_gnd_net_\,
            in3 => \N__41081\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41078\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46805\,
            in1 => \N__44092\,
            in2 => \_gnd_net_\,
            in3 => \N__41064\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44609\,
            in1 => \N__46945\,
            in2 => \N__45253\,
            in3 => \N__41148\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44088\,
            in1 => \N__46046\,
            in2 => \_gnd_net_\,
            in3 => \N__43650\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__44592\,
            in1 => \_gnd_net_\,
            in2 => \N__48159\,
            in3 => \N__44193\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__45258\,
            in1 => \N__44591\,
            in2 => \N__45428\,
            in3 => \N__46292\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44593\,
            in1 => \N__47991\,
            in2 => \_gnd_net_\,
            in3 => \N__41272\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47907\,
            in1 => \N__44594\,
            in2 => \_gnd_net_\,
            in3 => \N__44145\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__43611\,
            in1 => \N__44087\,
            in2 => \_gnd_net_\,
            in3 => \N__46344\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46558\,
            in2 => \N__44098\,
            in3 => \N__45368\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44590\,
            in1 => \N__45259\,
            in2 => \N__43886\,
            in3 => \N__45477\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__41208\,
            in1 => \N__44086\,
            in2 => \_gnd_net_\,
            in3 => \N__46412\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46343\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44610\,
            in1 => \N__46935\,
            in2 => \N__45288\,
            in3 => \N__41155\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46858\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46735\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46473\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46215\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46929\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48140\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46154\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46542\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46095\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48219\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46605\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47981\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47897\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48066\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001110"
        )
    port map (
            in0 => \N__41805\,
            in1 => \N__41587\,
            in2 => \N__41906\,
            in3 => \N__41432\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__41885\,
            in1 => \N__41861\,
            in2 => \N__41824\,
            in3 => \N__41588\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__41503\,
            in1 => \N__41441\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIPFL2M1_0_1\,
            ltout => \elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__42220\,
            in1 => \N__41414\,
            in2 => \N__41402\,
            in3 => \N__41399\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47864\,
            ce => \N__43368\,
            sr => \N__47284\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__42534\,
            in1 => \N__42296\,
            in2 => \N__42240\,
            in3 => \N__42691\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47864\,
            ce => \N__43368\,
            sr => \N__47284\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__42221\,
            in1 => \N__42661\,
            in2 => \N__42307\,
            in3 => \N__42536\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47864\,
            ce => \N__43368\,
            sr => \N__47284\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__42533\,
            in1 => \N__42295\,
            in2 => \N__42586\,
            in3 => \N__42223\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47864\,
            ce => \N__43368\,
            sr => \N__47284\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__42222\,
            in1 => \N__42535\,
            in2 => \N__42308\,
            in3 => \N__42377\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47864\,
            ce => \N__43368\,
            sr => \N__47284\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__42532\,
            in1 => \N__42294\,
            in2 => \_gnd_net_\,
            in3 => \N__42625\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47864\,
            ce => \N__43368\,
            sr => \N__47284\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__42530\,
            in1 => \N__42232\,
            in2 => \N__42587\,
            in3 => \N__42293\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47859\,
            ce => \N__42115\,
            sr => \N__47289\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__42291\,
            in1 => \N__42531\,
            in2 => \N__42241\,
            in3 => \N__42373\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47859\,
            ce => \N__42115\,
            sr => \N__47289\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__42331\,
            in1 => \N__42292\,
            in2 => \N__42242\,
            in3 => \N__42170\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47859\,
            ce => \N__42115\,
            sr => \N__47289\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIM28A1_0_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__43061\,
            in1 => \N__42971\,
            in2 => \_gnd_net_\,
            in3 => \N__43030\,
            lcout => \phase_controller_inst1.stoper_tr.running_1_sqmuxa\,
            ltout => \phase_controller_inst1.stoper_tr.running_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__43031\,
            in1 => \N__42979\,
            in2 => \N__42914\,
            in3 => \N__42911\,
            lcout => \phase_controller_inst1.stoper_tr.un1_start_latched2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42866\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42844\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42806\,
            in2 => \N__42800\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43333\,
            in1 => \N__42764\,
            in2 => \_gnd_net_\,
            in3 => \N__42752\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__47846\,
            ce => 'H',
            sr => \N__47295\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__43337\,
            in1 => \N__42749\,
            in2 => \N__42743\,
            in3 => \N__42728\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__47846\,
            ce => 'H',
            sr => \N__47295\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43334\,
            in1 => \N__42725\,
            in2 => \_gnd_net_\,
            in3 => \N__42713\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__47846\,
            ce => 'H',
            sr => \N__47295\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43338\,
            in1 => \N__42710\,
            in2 => \_gnd_net_\,
            in3 => \N__42698\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__47846\,
            ce => 'H',
            sr => \N__47295\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43335\,
            in1 => \N__43181\,
            in2 => \_gnd_net_\,
            in3 => \N__43169\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__47846\,
            ce => 'H',
            sr => \N__47295\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43339\,
            in1 => \N__43166\,
            in2 => \_gnd_net_\,
            in3 => \N__43154\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__47846\,
            ce => 'H',
            sr => \N__47295\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43336\,
            in1 => \N__43151\,
            in2 => \_gnd_net_\,
            in3 => \N__43139\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__47846\,
            ce => 'H',
            sr => \N__47295\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43372\,
            in1 => \N__43136\,
            in2 => \_gnd_net_\,
            in3 => \N__43124\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__47303\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43326\,
            in1 => \N__43121\,
            in2 => \_gnd_net_\,
            in3 => \N__43109\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__47303\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43369\,
            in1 => \N__43106\,
            in2 => \_gnd_net_\,
            in3 => \N__43094\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__47303\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43327\,
            in1 => \N__43091\,
            in2 => \_gnd_net_\,
            in3 => \N__43079\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__47303\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43370\,
            in1 => \N__43076\,
            in2 => \_gnd_net_\,
            in3 => \N__43064\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__47303\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43328\,
            in1 => \N__43448\,
            in2 => \_gnd_net_\,
            in3 => \N__43436\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__47303\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43371\,
            in1 => \N__43433\,
            in2 => \_gnd_net_\,
            in3 => \N__43421\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__47303\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43329\,
            in1 => \N__43418\,
            in2 => \_gnd_net_\,
            in3 => \N__43406\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__47303\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43330\,
            in1 => \N__43403\,
            in2 => \_gnd_net_\,
            in3 => \N__43391\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__47830\,
            ce => 'H',
            sr => \N__47307\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43332\,
            in1 => \N__43388\,
            in2 => \_gnd_net_\,
            in3 => \N__43376\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__47830\,
            ce => 'H',
            sr => \N__47307\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43331\,
            in1 => \N__43262\,
            in2 => \_gnd_net_\,
            in3 => \N__43265\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47830\,
            ce => 'H',
            sr => \N__47307\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44418\,
            in1 => \N__45837\,
            in2 => \N__45180\,
            in3 => \N__43250\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44075\,
            in1 => \N__46164\,
            in2 => \_gnd_net_\,
            in3 => \N__43497\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__45065\,
            in1 => \N__44456\,
            in2 => \N__43708\,
            in3 => \N__46111\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__43701\,
            in1 => \N__44076\,
            in2 => \_gnd_net_\,
            in3 => \N__46110\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__44457\,
            in1 => \N__46055\,
            in2 => \N__43663\,
            in3 => \N__45066\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44419\,
            in1 => \N__46351\,
            in2 => \N__45179\,
            in3 => \N__43612\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46298\,
            in1 => \N__44094\,
            in2 => \_gnd_net_\,
            in3 => \N__45417\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46227\,
            in1 => \N__44477\,
            in2 => \N__45264\,
            in3 => \N__43545\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44478\,
            in1 => \N__45215\,
            in2 => \N__43508\,
            in3 => \N__46165\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45899\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45603\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45211\,
            in1 => \N__44476\,
            in2 => \N__46490\,
            in3 => \N__43927\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45478\,
            in1 => \N__44093\,
            in2 => \_gnd_net_\,
            in3 => \N__43872\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45975\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__44463\,
            in1 => \N__43759\,
            in2 => \N__43811\,
            in3 => \N__43747\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45950\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47815\,
            ce => \N__47514\,
            sr => \N__47322\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43745\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__43748\,
            in1 => \N__44464\,
            in2 => \N__43763\,
            in3 => \N__43810\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__44078\,
            in1 => \N__43758\,
            in2 => \_gnd_net_\,
            in3 => \N__43746\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44465\,
            in2 => \_gnd_net_\,
            in3 => \N__44254\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__44255\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44579\,
            lcout => \current_shift_inst.un4_control_input_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44578\,
            in1 => \N__48237\,
            in2 => \_gnd_net_\,
            in3 => \N__45316\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45267\,
            in1 => \N__44576\,
            in2 => \N__48166\,
            in3 => \N__44197\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46419\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__45265\,
            in1 => \N__47914\,
            in2 => \N__44155\,
            in3 => \N__44577\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46293\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__46483\,
            in1 => \N__43931\,
            in2 => \N__45289\,
            in3 => \N__44573\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44099\,
            in1 => \N__46482\,
            in2 => \_gnd_net_\,
            in3 => \N__43923\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__45266\,
            in1 => \N__44575\,
            in2 => \N__46565\,
            in3 => \N__45366\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__44574\,
            in1 => \N__45271\,
            in2 => \N__45424\,
            in3 => \N__46294\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45470\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46050\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__44644\,
            in1 => \N__46557\,
            in2 => \N__45290\,
            in3 => \N__45367\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46682\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__48238\,
            in1 => \N__45315\,
            in2 => \N__45291\,
            in3 => \N__44645\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45669\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45529\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46018\,
            in2 => \N__45868\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__47797\,
            ce => \N__47513\,
            sr => \N__47332\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45946\,
            in2 => \N__45793\,
            in3 => \N__45872\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__47797\,
            ce => \N__47513\,
            sr => \N__47332\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45715\,
            in2 => \N__45869\,
            in3 => \N__45797\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__47797\,
            ce => \N__47513\,
            sr => \N__47332\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45646\,
            in2 => \N__45794\,
            in3 => \N__45722\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__47797\,
            ce => \N__47513\,
            sr => \N__47332\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45571\,
            in2 => \N__45719\,
            in3 => \N__45653\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__47797\,
            ce => \N__47513\,
            sr => \N__47332\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45511\,
            in2 => \N__45650\,
            in3 => \N__45578\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__47797\,
            ce => \N__47513\,
            sr => \N__47332\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46519\,
            in2 => \N__45575\,
            in3 => \N__45518\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__47797\,
            ce => \N__47513\,
            sr => \N__47332\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46453\,
            in2 => \N__45515\,
            in3 => \N__45449\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__47797\,
            ce => \N__47513\,
            sr => \N__47332\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46384\,
            in2 => \N__46523\,
            in3 => \N__46460\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__47792\,
            ce => \N__47512\,
            sr => \N__47334\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46318\,
            in2 => \N__46457\,
            in3 => \N__46391\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__47792\,
            ce => \N__47512\,
            sr => \N__47334\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46264\,
            in2 => \N__46388\,
            in3 => \N__46322\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__47792\,
            ce => \N__47512\,
            sr => \N__47334\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46319\,
            in2 => \N__46195\,
            in3 => \N__46271\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__47792\,
            ce => \N__47512\,
            sr => \N__47334\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46132\,
            in2 => \N__46268\,
            in3 => \N__46199\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__47792\,
            ce => \N__47512\,
            sr => \N__47334\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46075\,
            in2 => \N__46196\,
            in3 => \N__46136\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__47792\,
            ce => \N__47512\,
            sr => \N__47334\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46133\,
            in2 => \N__46981\,
            in3 => \N__46079\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__47792\,
            ce => \N__47512\,
            sr => \N__47334\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46076\,
            in2 => \N__46909\,
            in3 => \N__46022\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__47792\,
            ce => \N__47512\,
            sr => \N__47334\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46840\,
            in2 => \N__46982\,
            in3 => \N__46913\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__47787\,
            ce => \N__47511\,
            sr => \N__47340\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46771\,
            in2 => \N__46910\,
            in3 => \N__46847\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__47787\,
            ce => \N__47511\,
            sr => \N__47340\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46717\,
            in2 => \N__46844\,
            in3 => \N__46775\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__47787\,
            ce => \N__47511\,
            sr => \N__47340\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46772\,
            in2 => \N__46654\,
            in3 => \N__46724\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__47787\,
            ce => \N__47511\,
            sr => \N__47340\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46585\,
            in2 => \N__46721\,
            in3 => \N__46658\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__47787\,
            ce => \N__47511\,
            sr => \N__47340\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48262\,
            in2 => \N__46655\,
            in3 => \N__46589\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__47787\,
            ce => \N__47511\,
            sr => \N__47340\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46586\,
            in2 => \N__48202\,
            in3 => \N__46526\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__47787\,
            ce => \N__47511\,
            sr => \N__47340\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48263\,
            in2 => \N__48121\,
            in3 => \N__48206\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__47787\,
            ce => \N__47511\,
            sr => \N__47340\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48025\,
            in2 => \N__48203\,
            in3 => \N__48125\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_18_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__47783\,
            ce => \N__47510\,
            sr => \N__47351\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47938\,
            in2 => \N__48122\,
            in3 => \N__48050\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__47783\,
            ce => \N__47510\,
            sr => \N__47351\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48047\,
            in2 => \N__48029\,
            in3 => \N__47963\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__47783\,
            ce => \N__47510\,
            sr => \N__47351\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47960\,
            in2 => \N__47942\,
            in3 => \N__47879\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__47783\,
            ce => \N__47510\,
            sr => \N__47351\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47024\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
