// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 20 2025 00:15:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T12,
    s4_phy,
    rgb_g,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T12;
    output s4_phy;
    output rgb_g;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__21833;
    wire N__21832;
    wire N__21831;
    wire N__21822;
    wire N__21821;
    wire N__21820;
    wire N__21813;
    wire N__21812;
    wire N__21811;
    wire N__21804;
    wire N__21803;
    wire N__21802;
    wire N__21795;
    wire N__21794;
    wire N__21793;
    wire N__21786;
    wire N__21785;
    wire N__21784;
    wire N__21777;
    wire N__21776;
    wire N__21775;
    wire N__21768;
    wire N__21767;
    wire N__21766;
    wire N__21759;
    wire N__21758;
    wire N__21757;
    wire N__21750;
    wire N__21749;
    wire N__21748;
    wire N__21741;
    wire N__21740;
    wire N__21739;
    wire N__21732;
    wire N__21731;
    wire N__21730;
    wire N__21723;
    wire N__21722;
    wire N__21721;
    wire N__21714;
    wire N__21713;
    wire N__21712;
    wire N__21705;
    wire N__21704;
    wire N__21703;
    wire N__21686;
    wire N__21683;
    wire N__21682;
    wire N__21681;
    wire N__21680;
    wire N__21679;
    wire N__21678;
    wire N__21677;
    wire N__21676;
    wire N__21675;
    wire N__21672;
    wire N__21671;
    wire N__21670;
    wire N__21667;
    wire N__21666;
    wire N__21665;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21653;
    wire N__21646;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21628;
    wire N__21625;
    wire N__21620;
    wire N__21609;
    wire N__21606;
    wire N__21601;
    wire N__21596;
    wire N__21595;
    wire N__21594;
    wire N__21593;
    wire N__21592;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21560;
    wire N__21557;
    wire N__21556;
    wire N__21555;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21488;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21464;
    wire N__21463;
    wire N__21460;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21389;
    wire N__21388;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21377;
    wire N__21376;
    wire N__21375;
    wire N__21374;
    wire N__21373;
    wire N__21372;
    wire N__21371;
    wire N__21370;
    wire N__21369;
    wire N__21368;
    wire N__21367;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21350;
    wire N__21349;
    wire N__21348;
    wire N__21347;
    wire N__21346;
    wire N__21345;
    wire N__21344;
    wire N__21343;
    wire N__21340;
    wire N__21339;
    wire N__21338;
    wire N__21323;
    wire N__21318;
    wire N__21313;
    wire N__21312;
    wire N__21311;
    wire N__21300;
    wire N__21287;
    wire N__21282;
    wire N__21279;
    wire N__21274;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21250;
    wire N__21249;
    wire N__21248;
    wire N__21247;
    wire N__21246;
    wire N__21243;
    wire N__21232;
    wire N__21227;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21215;
    wire N__21214;
    wire N__21211;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21194;
    wire N__21193;
    wire N__21192;
    wire N__21191;
    wire N__21190;
    wire N__21189;
    wire N__21188;
    wire N__21187;
    wire N__21186;
    wire N__21185;
    wire N__21184;
    wire N__21183;
    wire N__21182;
    wire N__21181;
    wire N__21180;
    wire N__21179;
    wire N__21178;
    wire N__21177;
    wire N__21176;
    wire N__21175;
    wire N__21174;
    wire N__21173;
    wire N__21172;
    wire N__21171;
    wire N__21170;
    wire N__21169;
    wire N__21168;
    wire N__21167;
    wire N__21166;
    wire N__21165;
    wire N__21164;
    wire N__21163;
    wire N__21162;
    wire N__21161;
    wire N__21160;
    wire N__21159;
    wire N__21158;
    wire N__21157;
    wire N__21156;
    wire N__21155;
    wire N__21154;
    wire N__21153;
    wire N__21152;
    wire N__21151;
    wire N__21150;
    wire N__21149;
    wire N__21148;
    wire N__21147;
    wire N__21146;
    wire N__21145;
    wire N__21144;
    wire N__21143;
    wire N__21142;
    wire N__21141;
    wire N__21140;
    wire N__21139;
    wire N__21138;
    wire N__21137;
    wire N__21136;
    wire N__21135;
    wire N__21134;
    wire N__21133;
    wire N__21132;
    wire N__21131;
    wire N__21130;
    wire N__21129;
    wire N__21128;
    wire N__21127;
    wire N__21126;
    wire N__21125;
    wire N__21124;
    wire N__21123;
    wire N__21122;
    wire N__21121;
    wire N__21120;
    wire N__21119;
    wire N__21118;
    wire N__21117;
    wire N__21116;
    wire N__21115;
    wire N__21114;
    wire N__21113;
    wire N__21112;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21107;
    wire N__21106;
    wire N__21105;
    wire N__21104;
    wire N__21103;
    wire N__21102;
    wire N__21101;
    wire N__21100;
    wire N__21099;
    wire N__20906;
    wire N__20903;
    wire N__20902;
    wire N__20901;
    wire N__20900;
    wire N__20899;
    wire N__20898;
    wire N__20895;
    wire N__20894;
    wire N__20893;
    wire N__20892;
    wire N__20891;
    wire N__20890;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20846;
    wire N__20845;
    wire N__20844;
    wire N__20843;
    wire N__20840;
    wire N__20839;
    wire N__20838;
    wire N__20837;
    wire N__20836;
    wire N__20835;
    wire N__20834;
    wire N__20833;
    wire N__20832;
    wire N__20831;
    wire N__20830;
    wire N__20829;
    wire N__20828;
    wire N__20827;
    wire N__20826;
    wire N__20825;
    wire N__20824;
    wire N__20823;
    wire N__20822;
    wire N__20821;
    wire N__20820;
    wire N__20819;
    wire N__20818;
    wire N__20815;
    wire N__20814;
    wire N__20813;
    wire N__20812;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20808;
    wire N__20807;
    wire N__20806;
    wire N__20805;
    wire N__20804;
    wire N__20803;
    wire N__20802;
    wire N__20801;
    wire N__20800;
    wire N__20799;
    wire N__20798;
    wire N__20797;
    wire N__20796;
    wire N__20795;
    wire N__20794;
    wire N__20793;
    wire N__20792;
    wire N__20791;
    wire N__20790;
    wire N__20789;
    wire N__20788;
    wire N__20787;
    wire N__20786;
    wire N__20785;
    wire N__20784;
    wire N__20783;
    wire N__20782;
    wire N__20781;
    wire N__20780;
    wire N__20779;
    wire N__20778;
    wire N__20777;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20762;
    wire N__20761;
    wire N__20760;
    wire N__20759;
    wire N__20758;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20590;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20554;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20541;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20518;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20485;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20452;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20416;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20377;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20357;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20329;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20309;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20281;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20261;
    wire N__20260;
    wire N__20259;
    wire N__20258;
    wire N__20257;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20240;
    wire N__20237;
    wire N__20232;
    wire N__20229;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20213;
    wire N__20210;
    wire N__20209;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20189;
    wire N__20188;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20156;
    wire N__20153;
    wire N__20152;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20132;
    wire N__20131;
    wire N__20130;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20108;
    wire N__20105;
    wire N__20104;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20084;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20067;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20051;
    wire N__20048;
    wire N__20047;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20027;
    wire N__20026;
    wire N__20023;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20011;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19999;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19963;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19930;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19874;
    wire N__19871;
    wire N__19870;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19826;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19802;
    wire N__19801;
    wire N__19798;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19768;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19748;
    wire N__19745;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19723;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19703;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19682;
    wire N__19679;
    wire N__19678;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19658;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19637;
    wire N__19634;
    wire N__19633;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19613;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19586;
    wire N__19583;
    wire N__19582;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19562;
    wire N__19559;
    wire N__19558;
    wire N__19557;
    wire N__19556;
    wire N__19553;
    wire N__19548;
    wire N__19545;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19505;
    wire N__19504;
    wire N__19501;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19484;
    wire N__19481;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19463;
    wire N__19462;
    wire N__19461;
    wire N__19460;
    wire N__19459;
    wire N__19458;
    wire N__19457;
    wire N__19456;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19438;
    wire N__19437;
    wire N__19436;
    wire N__19435;
    wire N__19434;
    wire N__19433;
    wire N__19432;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19394;
    wire N__19393;
    wire N__19392;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19382;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19370;
    wire N__19353;
    wire N__19342;
    wire N__19339;
    wire N__19334;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19306;
    wire N__19305;
    wire N__19304;
    wire N__19303;
    wire N__19302;
    wire N__19301;
    wire N__19286;
    wire N__19285;
    wire N__19284;
    wire N__19283;
    wire N__19282;
    wire N__19281;
    wire N__19280;
    wire N__19279;
    wire N__19278;
    wire N__19277;
    wire N__19276;
    wire N__19275;
    wire N__19274;
    wire N__19273;
    wire N__19272;
    wire N__19269;
    wire N__19260;
    wire N__19257;
    wire N__19240;
    wire N__19239;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19227;
    wire N__19224;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19197;
    wire N__19184;
    wire N__19183;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19166;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19124;
    wire N__19121;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19097;
    wire N__19094;
    wire N__19093;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19073;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19049;
    wire N__19046;
    wire N__19045;
    wire N__19044;
    wire N__19041;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19025;
    wire N__19022;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19004;
    wire N__19001;
    wire N__19000;
    wire N__18999;
    wire N__18996;
    wire N__18993;
    wire N__18990;
    wire N__18987;
    wire N__18980;
    wire N__18977;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18969;
    wire N__18968;
    wire N__18963;
    wire N__18960;
    wire N__18957;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18937;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18920;
    wire N__18917;
    wire N__18912;
    wire N__18909;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18822;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18806;
    wire N__18805;
    wire N__18804;
    wire N__18803;
    wire N__18800;
    wire N__18795;
    wire N__18792;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18772;
    wire N__18769;
    wire N__18766;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18724;
    wire N__18723;
    wire N__18722;
    wire N__18721;
    wire N__18720;
    wire N__18719;
    wire N__18718;
    wire N__18717;
    wire N__18716;
    wire N__18715;
    wire N__18714;
    wire N__18713;
    wire N__18712;
    wire N__18711;
    wire N__18710;
    wire N__18709;
    wire N__18708;
    wire N__18707;
    wire N__18706;
    wire N__18705;
    wire N__18704;
    wire N__18703;
    wire N__18702;
    wire N__18701;
    wire N__18700;
    wire N__18699;
    wire N__18698;
    wire N__18697;
    wire N__18696;
    wire N__18687;
    wire N__18678;
    wire N__18669;
    wire N__18664;
    wire N__18655;
    wire N__18646;
    wire N__18637;
    wire N__18628;
    wire N__18621;
    wire N__18610;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18595;
    wire N__18594;
    wire N__18593;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18577;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18247;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18040;
    wire N__18039;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18024;
    wire N__18019;
    wire N__18016;
    wire N__18009;
    wire N__18006;
    wire N__18001;
    wire N__17996;
    wire N__17995;
    wire N__17992;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17978;
    wire N__17975;
    wire N__17974;
    wire N__17973;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17965;
    wire N__17964;
    wire N__17963;
    wire N__17962;
    wire N__17961;
    wire N__17960;
    wire N__17955;
    wire N__17950;
    wire N__17945;
    wire N__17936;
    wire N__17933;
    wire N__17926;
    wire N__17921;
    wire N__17920;
    wire N__17917;
    wire N__17916;
    wire N__17915;
    wire N__17914;
    wire N__17913;
    wire N__17908;
    wire N__17905;
    wire N__17902;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17884;
    wire N__17881;
    wire N__17880;
    wire N__17879;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17865;
    wire N__17858;
    wire N__17855;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17837;
    wire N__17834;
    wire N__17833;
    wire N__17832;
    wire N__17827;
    wire N__17826;
    wire N__17825;
    wire N__17822;
    wire N__17821;
    wire N__17820;
    wire N__17819;
    wire N__17818;
    wire N__17815;
    wire N__17806;
    wire N__17799;
    wire N__17798;
    wire N__17797;
    wire N__17796;
    wire N__17795;
    wire N__17794;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17745;
    wire N__17738;
    wire N__17735;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17722;
    wire N__17717;
    wire N__17716;
    wire N__17711;
    wire N__17710;
    wire N__17709;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17697;
    wire N__17690;
    wire N__17687;
    wire N__17686;
    wire N__17683;
    wire N__17682;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17660;
    wire N__17659;
    wire N__17658;
    wire N__17657;
    wire N__17656;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17638;
    wire N__17637;
    wire N__17636;
    wire N__17627;
    wire N__17626;
    wire N__17625;
    wire N__17624;
    wire N__17623;
    wire N__17622;
    wire N__17621;
    wire N__17620;
    wire N__17619;
    wire N__17618;
    wire N__17617;
    wire N__17614;
    wire N__17609;
    wire N__17600;
    wire N__17591;
    wire N__17590;
    wire N__17589;
    wire N__17588;
    wire N__17587;
    wire N__17578;
    wire N__17577;
    wire N__17576;
    wire N__17575;
    wire N__17574;
    wire N__17573;
    wire N__17572;
    wire N__17571;
    wire N__17570;
    wire N__17561;
    wire N__17558;
    wire N__17549;
    wire N__17540;
    wire N__17539;
    wire N__17538;
    wire N__17537;
    wire N__17536;
    wire N__17533;
    wire N__17526;
    wire N__17517;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17501;
    wire N__17500;
    wire N__17499;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17453;
    wire N__17452;
    wire N__17451;
    wire N__17448;
    wire N__17445;
    wire N__17442;
    wire N__17439;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17421;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17407;
    wire N__17404;
    wire N__17401;
    wire N__17400;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17370;
    wire N__17363;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17345;
    wire N__17342;
    wire N__17337;
    wire N__17334;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17313;
    wire N__17310;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17292;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17265;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17243;
    wire N__17242;
    wire N__17239;
    wire N__17238;
    wire N__17235;
    wire N__17234;
    wire N__17229;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17185;
    wire N__17184;
    wire N__17183;
    wire N__17180;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17146;
    wire N__17145;
    wire N__17142;
    wire N__17137;
    wire N__17132;
    wire N__17129;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17104;
    wire N__17103;
    wire N__17100;
    wire N__17095;
    wire N__17090;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17044;
    wire N__17041;
    wire N__17040;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16990;
    wire N__16985;
    wire N__16984;
    wire N__16983;
    wire N__16982;
    wire N__16981;
    wire N__16980;
    wire N__16977;
    wire N__16976;
    wire N__16975;
    wire N__16974;
    wire N__16971;
    wire N__16968;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16934;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16926;
    wire N__16925;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16900;
    wire N__16897;
    wire N__16892;
    wire N__16891;
    wire N__16888;
    wire N__16887;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16855;
    wire N__16850;
    wire N__16847;
    wire N__16846;
    wire N__16843;
    wire N__16840;
    wire N__16837;
    wire N__16836;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16792;
    wire N__16791;
    wire N__16790;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16776;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16743;
    wire N__16740;
    wire N__16737;
    wire N__16734;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16720;
    wire N__16719;
    wire N__16718;
    wire N__16717;
    wire N__16716;
    wire N__16715;
    wire N__16714;
    wire N__16713;
    wire N__16712;
    wire N__16711;
    wire N__16700;
    wire N__16697;
    wire N__16686;
    wire N__16685;
    wire N__16684;
    wire N__16683;
    wire N__16682;
    wire N__16681;
    wire N__16680;
    wire N__16679;
    wire N__16678;
    wire N__16677;
    wire N__16676;
    wire N__16675;
    wire N__16672;
    wire N__16667;
    wire N__16656;
    wire N__16643;
    wire N__16642;
    wire N__16639;
    wire N__16632;
    wire N__16629;
    wire N__16622;
    wire N__16621;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16610;
    wire N__16609;
    wire N__16608;
    wire N__16607;
    wire N__16606;
    wire N__16605;
    wire N__16604;
    wire N__16603;
    wire N__16602;
    wire N__16601;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16580;
    wire N__16579;
    wire N__16576;
    wire N__16567;
    wire N__16566;
    wire N__16565;
    wire N__16564;
    wire N__16563;
    wire N__16562;
    wire N__16559;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16531;
    wire N__16528;
    wire N__16521;
    wire N__16514;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16469;
    wire N__16468;
    wire N__16467;
    wire N__16464;
    wire N__16461;
    wire N__16458;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16441;
    wire N__16440;
    wire N__16439;
    wire N__16438;
    wire N__16437;
    wire N__16436;
    wire N__16435;
    wire N__16434;
    wire N__16431;
    wire N__16430;
    wire N__16429;
    wire N__16428;
    wire N__16425;
    wire N__16422;
    wire N__16419;
    wire N__16416;
    wire N__16415;
    wire N__16414;
    wire N__16413;
    wire N__16412;
    wire N__16401;
    wire N__16400;
    wire N__16399;
    wire N__16398;
    wire N__16393;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16373;
    wire N__16372;
    wire N__16371;
    wire N__16370;
    wire N__16367;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16356;
    wire N__16355;
    wire N__16352;
    wire N__16347;
    wire N__16330;
    wire N__16329;
    wire N__16326;
    wire N__16315;
    wire N__16310;
    wire N__16307;
    wire N__16298;
    wire N__16295;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16285;
    wire N__16284;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16272;
    wire N__16265;
    wire N__16262;
    wire N__16261;
    wire N__16260;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16232;
    wire N__16229;
    wire N__16228;
    wire N__16227;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16215;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16199;
    wire N__16196;
    wire N__16195;
    wire N__16194;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16176;
    wire N__16171;
    wire N__16166;
    wire N__16165;
    wire N__16162;
    wire N__16161;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16149;
    wire N__16146;
    wire N__16141;
    wire N__16136;
    wire N__16133;
    wire N__16132;
    wire N__16127;
    wire N__16124;
    wire N__16123;
    wire N__16122;
    wire N__16119;
    wire N__16114;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16102;
    wire N__16101;
    wire N__16098;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16084;
    wire N__16081;
    wire N__16076;
    wire N__16071;
    wire N__16064;
    wire N__16063;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16053;
    wire N__16052;
    wire N__16051;
    wire N__16048;
    wire N__16043;
    wire N__16038;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16015;
    wire N__16012;
    wire N__16011;
    wire N__16006;
    wire N__16005;
    wire N__16002;
    wire N__15999;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15973;
    wire N__15972;
    wire N__15969;
    wire N__15966;
    wire N__15963;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15938;
    wire N__15937;
    wire N__15936;
    wire N__15935;
    wire N__15930;
    wire N__15927;
    wire N__15926;
    wire N__15923;
    wire N__15922;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15908;
    wire N__15899;
    wire N__15898;
    wire N__15897;
    wire N__15894;
    wire N__15891;
    wire N__15890;
    wire N__15889;
    wire N__15888;
    wire N__15887;
    wire N__15886;
    wire N__15885;
    wire N__15884;
    wire N__15883;
    wire N__15882;
    wire N__15879;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15855;
    wire N__15854;
    wire N__15853;
    wire N__15852;
    wire N__15851;
    wire N__15850;
    wire N__15849;
    wire N__15846;
    wire N__15843;
    wire N__15840;
    wire N__15835;
    wire N__15834;
    wire N__15833;
    wire N__15832;
    wire N__15831;
    wire N__15830;
    wire N__15829;
    wire N__15828;
    wire N__15827;
    wire N__15824;
    wire N__15817;
    wire N__15810;
    wire N__15807;
    wire N__15800;
    wire N__15783;
    wire N__15778;
    wire N__15767;
    wire N__15764;
    wire N__15763;
    wire N__15762;
    wire N__15761;
    wire N__15756;
    wire N__15753;
    wire N__15750;
    wire N__15743;
    wire N__15742;
    wire N__15741;
    wire N__15740;
    wire N__15739;
    wire N__15738;
    wire N__15737;
    wire N__15736;
    wire N__15735;
    wire N__15734;
    wire N__15733;
    wire N__15732;
    wire N__15731;
    wire N__15730;
    wire N__15729;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15715;
    wire N__15714;
    wire N__15713;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15687;
    wire N__15686;
    wire N__15669;
    wire N__15666;
    wire N__15657;
    wire N__15648;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15626;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15610;
    wire N__15607;
    wire N__15604;
    wire N__15593;
    wire N__15592;
    wire N__15591;
    wire N__15590;
    wire N__15589;
    wire N__15588;
    wire N__15587;
    wire N__15586;
    wire N__15569;
    wire N__15568;
    wire N__15567;
    wire N__15566;
    wire N__15563;
    wire N__15562;
    wire N__15561;
    wire N__15560;
    wire N__15559;
    wire N__15558;
    wire N__15557;
    wire N__15556;
    wire N__15555;
    wire N__15554;
    wire N__15553;
    wire N__15552;
    wire N__15551;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15529;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15481;
    wire N__15478;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15461;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15433;
    wire N__15432;
    wire N__15425;
    wire N__15422;
    wire N__15421;
    wire N__15420;
    wire N__15419;
    wire N__15416;
    wire N__15409;
    wire N__15404;
    wire N__15401;
    wire N__15400;
    wire N__15397;
    wire N__15394;
    wire N__15389;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15365;
    wire N__15364;
    wire N__15363;
    wire N__15362;
    wire N__15361;
    wire N__15356;
    wire N__15349;
    wire N__15344;
    wire N__15343;
    wire N__15340;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15325;
    wire N__15322;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15305;
    wire N__15302;
    wire N__15301;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15289;
    wire N__15284;
    wire N__15283;
    wire N__15282;
    wire N__15281;
    wire N__15280;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15272;
    wire N__15269;
    wire N__15264;
    wire N__15259;
    wire N__15252;
    wire N__15245;
    wire N__15244;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15215;
    wire N__15214;
    wire N__15211;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15196;
    wire N__15191;
    wire N__15190;
    wire N__15189;
    wire N__15186;
    wire N__15181;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15142;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15116;
    wire N__15113;
    wire N__15112;
    wire N__15111;
    wire N__15108;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15071;
    wire N__15068;
    wire N__15067;
    wire N__15066;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15056;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15042;
    wire N__15037;
    wire N__15032;
    wire N__15029;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15021;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15009;
    wire N__15004;
    wire N__15001;
    wire N__14996;
    wire N__14995;
    wire N__14992;
    wire N__14991;
    wire N__14990;
    wire N__14989;
    wire N__14988;
    wire N__14987;
    wire N__14984;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14970;
    wire N__14963;
    wire N__14960;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14948;
    wire N__14947;
    wire N__14946;
    wire N__14945;
    wire N__14942;
    wire N__14935;
    wire N__14928;
    wire N__14925;
    wire N__14918;
    wire N__14915;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14907;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14895;
    wire N__14892;
    wire N__14887;
    wire N__14882;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14862;
    wire N__14857;
    wire N__14854;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14842;
    wire N__14841;
    wire N__14838;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14814;
    wire N__14807;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14410;
    wire N__14407;
    wire N__14404;
    wire N__14399;
    wire N__14398;
    wire N__14397;
    wire N__14394;
    wire N__14391;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14369;
    wire N__14366;
    wire N__14365;
    wire N__14364;
    wire N__14361;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14345;
    wire N__14342;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14330;
    wire N__14327;
    wire N__14326;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14303;
    wire N__14302;
    wire N__14301;
    wire N__14300;
    wire N__14299;
    wire N__14296;
    wire N__14287;
    wire N__14284;
    wire N__14283;
    wire N__14280;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14258;
    wire N__14257;
    wire N__14256;
    wire N__14255;
    wire N__14254;
    wire N__14253;
    wire N__14252;
    wire N__14251;
    wire N__14242;
    wire N__14237;
    wire N__14232;
    wire N__14225;
    wire N__14224;
    wire N__14223;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14215;
    wire N__14212;
    wire N__14211;
    wire N__14210;
    wire N__14201;
    wire N__14196;
    wire N__14193;
    wire N__14186;
    wire N__14183;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14171;
    wire N__14168;
    wire N__14167;
    wire N__14166;
    wire N__14163;
    wire N__14158;
    wire N__14153;
    wire N__14152;
    wire N__14151;
    wire N__14148;
    wire N__14143;
    wire N__14138;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14130;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14116;
    wire N__14115;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14103;
    wire N__14100;
    wire N__14095;
    wire N__14090;
    wire N__14087;
    wire N__14086;
    wire N__14083;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14045;
    wire N__14042;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14027;
    wire N__14026;
    wire N__14025;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13882;
    wire N__13881;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13869;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13852;
    wire N__13851;
    wire N__13850;
    wire N__13845;
    wire N__13842;
    wire N__13839;
    wire N__13834;
    wire N__13831;
    wire N__13828;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13805;
    wire N__13802;
    wire N__13799;
    wire N__13798;
    wire N__13795;
    wire N__13794;
    wire N__13793;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13769;
    wire N__13760;
    wire N__13757;
    wire N__13754;
    wire N__13753;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13727;
    wire N__13726;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13718;
    wire N__13715;
    wire N__13714;
    wire N__13713;
    wire N__13712;
    wire N__13709;
    wire N__13704;
    wire N__13701;
    wire N__13698;
    wire N__13695;
    wire N__13692;
    wire N__13691;
    wire N__13688;
    wire N__13687;
    wire N__13684;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13656;
    wire N__13649;
    wire N__13648;
    wire N__13645;
    wire N__13642;
    wire N__13641;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13613;
    wire N__13612;
    wire N__13611;
    wire N__13608;
    wire N__13605;
    wire N__13602;
    wire N__13601;
    wire N__13598;
    wire N__13593;
    wire N__13590;
    wire N__13583;
    wire N__13580;
    wire N__13579;
    wire N__13576;
    wire N__13575;
    wire N__13572;
    wire N__13569;
    wire N__13566;
    wire N__13563;
    wire N__13558;
    wire N__13557;
    wire N__13552;
    wire N__13549;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13537;
    wire N__13534;
    wire N__13531;
    wire N__13530;
    wire N__13527;
    wire N__13524;
    wire N__13521;
    wire N__13518;
    wire N__13513;
    wire N__13508;
    wire N__13505;
    wire N__13504;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13472;
    wire N__13469;
    wire N__13468;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13458;
    wire N__13457;
    wire N__13456;
    wire N__13453;
    wire N__13450;
    wire N__13447;
    wire N__13444;
    wire N__13441;
    wire N__13430;
    wire N__13427;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13419;
    wire N__13418;
    wire N__13413;
    wire N__13408;
    wire N__13405;
    wire N__13402;
    wire N__13397;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13385;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13375;
    wire N__13372;
    wire N__13369;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13354;
    wire N__13351;
    wire N__13348;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13288;
    wire N__13287;
    wire N__13286;
    wire N__13285;
    wire N__13284;
    wire N__13283;
    wire N__13282;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13274;
    wire N__13273;
    wire N__13272;
    wire N__13271;
    wire N__13256;
    wire N__13255;
    wire N__13254;
    wire N__13253;
    wire N__13252;
    wire N__13251;
    wire N__13250;
    wire N__13249;
    wire N__13248;
    wire N__13245;
    wire N__13242;
    wire N__13239;
    wire N__13236;
    wire N__13233;
    wire N__13230;
    wire N__13229;
    wire N__13228;
    wire N__13227;
    wire N__13226;
    wire N__13225;
    wire N__13222;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13178;
    wire N__13163;
    wire N__13162;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13152;
    wire N__13145;
    wire N__13142;
    wire N__13141;
    wire N__13140;
    wire N__13139;
    wire N__13138;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13122;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13060;
    wire N__13057;
    wire N__13054;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13039;
    wire N__13036;
    wire N__13033;
    wire N__13028;
    wire N__13025;
    wire N__13022;
    wire N__13019;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12901;
    wire N__12898;
    wire N__12895;
    wire N__12892;
    wire N__12889;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12832;
    wire N__12829;
    wire N__12826;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12802;
    wire N__12799;
    wire N__12796;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12772;
    wire N__12769;
    wire N__12766;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12697;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12679;
    wire N__12676;
    wire N__12671;
    wire N__12668;
    wire N__12667;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12651;
    wire N__12644;
    wire N__12643;
    wire N__12640;
    wire N__12637;
    wire N__12632;
    wire N__12631;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12623;
    wire N__12620;
    wire N__12615;
    wire N__12612;
    wire N__12611;
    wire N__12608;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12508;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12487;
    wire N__12484;
    wire N__12481;
    wire N__12476;
    wire N__12473;
    wire N__12472;
    wire N__12469;
    wire N__12466;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12451;
    wire N__12448;
    wire N__12445;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12356;
    wire N__12353;
    wire N__12350;
    wire N__12347;
    wire N__12344;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12334;
    wire N__12329;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12280;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12188;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12173;
    wire N__12170;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12127;
    wire N__12124;
    wire N__12121;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12031;
    wire N__12030;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12016;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11994;
    wire N__11991;
    wire N__11984;
    wire N__11981;
    wire N__11980;
    wire N__11977;
    wire N__11974;
    wire N__11973;
    wire N__11968;
    wire N__11965;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11900;
    wire N__11899;
    wire N__11898;
    wire N__11897;
    wire N__11894;
    wire N__11893;
    wire N__11892;
    wire N__11891;
    wire N__11890;
    wire N__11883;
    wire N__11878;
    wire N__11877;
    wire N__11876;
    wire N__11875;
    wire N__11874;
    wire N__11873;
    wire N__11872;
    wire N__11869;
    wire N__11864;
    wire N__11861;
    wire N__11858;
    wire N__11847;
    wire N__11844;
    wire N__11843;
    wire N__11842;
    wire N__11841;
    wire N__11840;
    wire N__11839;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11825;
    wire N__11818;
    wire N__11811;
    wire N__11808;
    wire N__11803;
    wire N__11800;
    wire N__11789;
    wire N__11788;
    wire N__11787;
    wire N__11786;
    wire N__11785;
    wire N__11784;
    wire N__11783;
    wire N__11782;
    wire N__11781;
    wire N__11778;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11770;
    wire N__11767;
    wire N__11764;
    wire N__11763;
    wire N__11762;
    wire N__11761;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11751;
    wire N__11750;
    wire N__11749;
    wire N__11748;
    wire N__11747;
    wire N__11746;
    wire N__11745;
    wire N__11742;
    wire N__11735;
    wire N__11724;
    wire N__11717;
    wire N__11708;
    wire N__11707;
    wire N__11706;
    wire N__11703;
    wire N__11702;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11689;
    wire N__11686;
    wire N__11683;
    wire N__11676;
    wire N__11675;
    wire N__11674;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11658;
    wire N__11651;
    wire N__11644;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11618;
    wire N__11617;
    wire N__11616;
    wire N__11615;
    wire N__11614;
    wire N__11613;
    wire N__11612;
    wire N__11611;
    wire N__11610;
    wire N__11609;
    wire N__11602;
    wire N__11591;
    wire N__11586;
    wire N__11585;
    wire N__11584;
    wire N__11583;
    wire N__11582;
    wire N__11581;
    wire N__11580;
    wire N__11579;
    wire N__11578;
    wire N__11577;
    wire N__11576;
    wire N__11575;
    wire N__11572;
    wire N__11567;
    wire N__11560;
    wire N__11551;
    wire N__11542;
    wire N__11541;
    wire N__11540;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11476;
    wire N__11475;
    wire N__11474;
    wire N__11473;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11469;
    wire N__11468;
    wire N__11467;
    wire N__11466;
    wire N__11465;
    wire N__11464;
    wire N__11463;
    wire N__11462;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11458;
    wire N__11441;
    wire N__11430;
    wire N__11429;
    wire N__11428;
    wire N__11427;
    wire N__11426;
    wire N__11411;
    wire N__11406;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11387;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11365;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11361;
    wire N__11360;
    wire N__11359;
    wire N__11358;
    wire N__11357;
    wire N__11356;
    wire N__11353;
    wire N__11352;
    wire N__11351;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11337;
    wire N__11334;
    wire N__11333;
    wire N__11332;
    wire N__11331;
    wire N__11326;
    wire N__11325;
    wire N__11324;
    wire N__11323;
    wire N__11322;
    wire N__11319;
    wire N__11316;
    wire N__11313;
    wire N__11312;
    wire N__11309;
    wire N__11294;
    wire N__11283;
    wire N__11280;
    wire N__11263;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11239;
    wire N__11236;
    wire N__11231;
    wire N__11230;
    wire N__11227;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11215;
    wire N__11210;
    wire N__11207;
    wire N__11206;
    wire N__11203;
    wire N__11202;
    wire N__11199;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11187;
    wire N__11182;
    wire N__11181;
    wire N__11176;
    wire N__11173;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11053;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11038;
    wire N__11033;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11014;
    wire N__11009;
    wire N__11006;
    wire N__11005;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10988;
    wire N__10985;
    wire N__10984;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10967;
    wire N__10964;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10952;
    wire N__10951;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10941;
    wire N__10936;
    wire N__10931;
    wire N__10928;
    wire N__10927;
    wire N__10924;
    wire N__10921;
    wire N__10916;
    wire N__10915;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10900;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10885;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10858;
    wire N__10857;
    wire N__10854;
    wire N__10849;
    wire N__10844;
    wire N__10841;
    wire N__10840;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10825;
    wire N__10820;
    wire N__10817;
    wire N__10816;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10801;
    wire N__10796;
    wire N__10793;
    wire N__10792;
    wire N__10791;
    wire N__10788;
    wire N__10785;
    wire N__10782;
    wire N__10775;
    wire N__10772;
    wire N__10771;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10761;
    wire N__10754;
    wire N__10751;
    wire N__10750;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10735;
    wire N__10730;
    wire N__10727;
    wire N__10726;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10711;
    wire N__10706;
    wire N__10703;
    wire N__10702;
    wire N__10701;
    wire N__10698;
    wire N__10693;
    wire N__10688;
    wire N__10685;
    wire N__10684;
    wire N__10683;
    wire N__10680;
    wire N__10675;
    wire N__10670;
    wire N__10667;
    wire N__10666;
    wire N__10665;
    wire N__10662;
    wire N__10657;
    wire N__10652;
    wire N__10649;
    wire N__10648;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10638;
    wire N__10633;
    wire N__10628;
    wire N__10625;
    wire N__10624;
    wire N__10623;
    wire N__10620;
    wire N__10617;
    wire N__10614;
    wire N__10609;
    wire N__10604;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10583;
    wire N__10580;
    wire N__10579;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10562;
    wire N__10559;
    wire N__10558;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10543;
    wire N__10538;
    wire N__10535;
    wire N__10534;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10519;
    wire N__10514;
    wire N__10511;
    wire N__10510;
    wire N__10509;
    wire N__10506;
    wire N__10501;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10489;
    wire N__10488;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10472;
    wire N__10471;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10454;
    wire N__10451;
    wire N__10450;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10435;
    wire N__10430;
    wire N__10427;
    wire N__10426;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10411;
    wire N__10406;
    wire N__10403;
    wire N__10402;
    wire N__10401;
    wire N__10398;
    wire N__10393;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10159;
    wire N__10158;
    wire N__10157;
    wire N__10152;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9865;
    wire N__9864;
    wire N__9863;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9847;
    wire N__9842;
    wire N__9839;
    wire N__9838;
    wire N__9835;
    wire N__9832;
    wire N__9827;
    wire N__9824;
    wire N__9823;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9771;
    wire N__9768;
    wire N__9765;
    wire N__9762;
    wire N__9755;
    wire N__9752;
    wire N__9751;
    wire N__9750;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9685;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9658;
    wire N__9657;
    wire N__9652;
    wire N__9649;
    wire N__9644;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9636;
    wire N__9631;
    wire N__9628;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9583;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9575;
    wire N__9572;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9549;
    wire N__9546;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9418;
    wire N__9417;
    wire N__9416;
    wire N__9415;
    wire N__9414;
    wire N__9411;
    wire N__9400;
    wire N__9395;
    wire N__9392;
    wire N__9391;
    wire N__9390;
    wire N__9387;
    wire N__9384;
    wire N__9381;
    wire N__9374;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8953;
    wire N__8952;
    wire N__8951;
    wire N__8950;
    wire N__8949;
    wire N__8948;
    wire N__8947;
    wire N__8946;
    wire N__8945;
    wire N__8942;
    wire N__8941;
    wire N__8940;
    wire N__8939;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8928;
    wire N__8927;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8913;
    wire N__8912;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8904;
    wire N__8903;
    wire N__8902;
    wire N__8899;
    wire N__8884;
    wire N__8881;
    wire N__8876;
    wire N__8861;
    wire N__8850;
    wire N__8847;
    wire N__8840;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8818;
    wire N__8817;
    wire N__8816;
    wire N__8813;
    wire N__8812;
    wire N__8811;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8800;
    wire N__8799;
    wire N__8798;
    wire N__8797;
    wire N__8796;
    wire N__8795;
    wire N__8794;
    wire N__8793;
    wire N__8792;
    wire N__8791;
    wire N__8790;
    wire N__8789;
    wire N__8786;
    wire N__8781;
    wire N__8780;
    wire N__8779;
    wire N__8778;
    wire N__8777;
    wire N__8774;
    wire N__8773;
    wire N__8766;
    wire N__8763;
    wire N__8762;
    wire N__8761;
    wire N__8746;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8718;
    wire N__8713;
    wire N__8708;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8683;
    wire N__8682;
    wire N__8681;
    wire N__8680;
    wire N__8679;
    wire N__8678;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8671;
    wire N__8670;
    wire N__8669;
    wire N__8668;
    wire N__8667;
    wire N__8666;
    wire N__8665;
    wire N__8650;
    wire N__8649;
    wire N__8648;
    wire N__8633;
    wire N__8622;
    wire N__8621;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8608;
    wire N__8603;
    wire N__8598;
    wire N__8585;
    wire N__8584;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8374;
    wire N__8373;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_18_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_1_19_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_1_20_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire N_39_i_i;
    wire CONSTANT_ONE_NET;
    wire rgb_drv_RNOZ0;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUSZ0Z53 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.stoper_tr.N_60 ;
    wire \phase_controller_slave.start_timer_trZ0 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_1 ;
    wire bfn_3_18_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_9 ;
    wire bfn_3_19_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_17 ;
    wire bfn_3_20_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.tr_time_passed ;
    wire \phase_controller_slave.stateZ0Z_0 ;
    wire \phase_controller_slave.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ1Z_6 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1 ;
    wire il_max_comp2_c;
    wire il_min_comp2_c;
    wire il_min_comp2_D1;
    wire il_max_comp2_D1;
    wire \phase_controller_slave.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_slave.start_timer_hc_RNOZ0Z_0 ;
    wire il_min_comp2_D2;
    wire \phase_controller_slave.stateZ0Z_2 ;
    wire il_max_comp2_D2;
    wire \phase_controller_slave.stoper_hc.N_60 ;
    wire \phase_controller_slave.hc_time_passed ;
    wire \phase_controller_slave.state_RNIVDE2Z0Z_0 ;
    wire \phase_controller_slave.stateZ0Z_4 ;
    wire \phase_controller_slave.state_RNO_0Z0Z_3 ;
    wire shift_flag_start;
    wire \phase_controller_slave.stateZ0Z_1 ;
    wire s4_phy_c;
    wire bfn_7_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_7_14_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_7_15_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_7_16_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire bfn_7_17_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire bfn_7_18_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire bfn_7_19_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un1_startlt8_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_startlto5Z0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.un2_startlto6Z0Z_0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un2_startlt19_0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_start ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_7_23_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ1Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_7_24_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_7_25_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire il_max_comp1_c;
    wire \delay_measurement_inst.delay_hc_timer.N_105_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_8_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_8_14_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_8_15_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_8_16_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_178_i_g ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DKZ0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \phase_controller_slave.start_timer_hcZ0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_startlto9_cZ0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_startlto13 ;
    wire \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un3_start ;
    wire \phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_startlt15 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire bfn_8_25_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire bfn_8_26_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire bfn_8_27_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \delay_measurement_inst.delay_tr_timer.N_180_i ;
    wire il_min_comp1_c;
    wire \delay_measurement_inst.delay_hc_timer.N_101 ;
    wire \delay_measurement_inst.delay_hc_timer.N_81_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_5 ;
    wire \delay_measurement_inst.delay_hc_timer.N_105 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_0 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_9_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire measured_delay_tr_8;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_7_9 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_6_9_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_0_9 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_1 ;
    wire bfn_9_17_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_9 ;
    wire bfn_9_18_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_17 ;
    wire bfn_9_19_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire il_min_comp1_D1;
    wire measured_delay_tr_15;
    wire measured_delay_tr_6;
    wire measured_delay_tr_12;
    wire measured_delay_tr_14;
    wire measured_delay_tr_1;
    wire measured_delay_tr_17;
    wire measured_delay_tr_9;
    wire measured_delay_tr_5;
    wire \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_5_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_9_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_160_cascade_ ;
    wire \delay_measurement_inst.tr_state_RNIVV8GZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_reset_i_0 ;
    wire \phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_2 ;
    wire measured_delay_tr_7;
    wire measured_delay_tr_16;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stateZ0Z_3 ;
    wire s3_phy_c;
    wire \delay_measurement_inst.N_54_cascade_ ;
    wire \delay_measurement_inst.tr_syncZ0Z_1 ;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire \delay_measurement_inst.tr_prevZ0 ;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_hc_14 ;
    wire \delay_measurement_inst.elapsed_time_hc_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.N_32 ;
    wire \delay_measurement_inst.N_54_i ;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.N_109 ;
    wire \delay_measurement_inst.N_45 ;
    wire \delay_measurement_inst.N_107 ;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_10_15_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_10_16_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire bfn_10_17_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.stoper_state_RNI10KLZ0Z_1 ;
    wire measured_delay_tr_3;
    wire measured_delay_tr_18;
    wire measured_delay_tr_4;
    wire \delay_measurement_inst.N_129 ;
    wire \delay_measurement_inst.N_172 ;
    wire measured_delay_tr_2;
    wire measured_delay_tr_10;
    wire measured_delay_tr_11;
    wire measured_delay_tr_13;
    wire \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_6 ;
    wire \delay_measurement_inst.N_132 ;
    wire \delay_measurement_inst.N_139 ;
    wire \delay_measurement_inst.N_134_i ;
    wire \delay_measurement_inst.N_201_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_167 ;
    wire \delay_measurement_inst.N_170 ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.T01_0_sqmuxa ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire T12_c;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.N_60 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_181_i ;
    wire \delay_measurement_inst.hc_prevZ0 ;
    wire \delay_measurement_inst.hc_syncZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.N_81 ;
    wire \delay_measurement_inst.N_54 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt8_cascade_ ;
    wire measured_delay_hc_8;
    wire measured_delay_hc_7;
    wire \phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto13 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8_cascade_ ;
    wire measured_delay_hc_1;
    wire \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_2 ;
    wire measured_delay_hc_5;
    wire measured_delay_hc_16;
    wire measured_delay_hc_19;
    wire measured_delay_hc_17;
    wire measured_delay_hc_18;
    wire \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_start ;
    wire measured_delay_hc_6;
    wire \phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire measured_delay_hc_9;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire measured_delay_hc_13;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt15 ;
    wire \phase_controller_inst1.stoper_hc.un3_start ;
    wire measured_delay_hc_10;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire measured_delay_hc_14;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.N_201 ;
    wire measured_delay_tr_19;
    wire \delay_measurement_inst.N_134_i_0 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_7_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_4 ;
    wire \delay_measurement_inst.delay_tr_timer.N_127 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_6_9 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_0_9 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire delay_hc_d2;
    wire \delay_measurement_inst.hc_syncZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.elapsed_time_hc_15 ;
    wire \delay_measurement_inst.N_84 ;
    wire \delay_measurement_inst.N_40 ;
    wire measured_delay_hc_15;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire \delay_measurement_inst.N_48 ;
    wire \delay_measurement_inst.N_54_i_0 ;
    wire \delay_measurement_inst.N_32_g ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.N_179_i_g ;
    wire measured_delay_hc_2;
    wire \phase_controller_inst1.stoper_hc.un2_startlto6Z0Z_0 ;
    wire measured_delay_hc_3;
    wire measured_delay_hc_4;
    wire \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_4 ;
    wire measured_delay_hc_12;
    wire \phase_controller_inst1.stoper_hc.un2_startlt19_0_cascade_ ;
    wire measured_delay_hc_11;
    wire \phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9 ;
    wire il_max_comp1_D1;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire bfn_12_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire bfn_12_16_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire bfn_12_17_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire bfn_12_18_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_12_19_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_12_20_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_12_21_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_181_i_g ;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.N_108 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \phase_controller_inst1.stateZ0Z_3 ;
    wire s1_phy_c;
    wire \pll_inst.red_c_i ;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire \delay_measurement_inst.tr_syncZ0Z_0 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_178_i ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.N_112 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire bfn_13_19_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire bfn_13_20_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.elapsed_time_tr_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.elapsed_time_tr_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire bfn_13_21_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_13_22_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.N_180_i_g ;
    wire start_stop_c;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \phase_controller_inst1.N_110 ;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire T23_c;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.N_60 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire _gnd_net_;
    wire clk_100mhz;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__17066),
            .RESETB(N__18890),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__21831),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__21833),
            .DIN(N__21832),
            .DOUT(N__21831),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__21833),
            .PADOUT(N__21832),
            .PADIN(N__21831),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__21822),
            .DIN(N__21821),
            .DOUT(N__21820),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__21822),
            .PADOUT(N__21821),
            .PADIN(N__21820),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__21813),
            .DIN(N__21812),
            .DOUT(N__21811),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__21813),
            .PADOUT(N__21812),
            .PADIN(N__21811),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18902),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__21804),
            .DIN(N__21803),
            .DOUT(N__21802),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__21804),
            .PADOUT(N__21803),
            .PADIN(N__21802),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9728),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__21795),
            .DIN(N__21794),
            .DOUT(N__21793),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__21795),
            .PADOUT(N__21794),
            .PADIN(N__21793),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__21786),
            .DIN(N__21785),
            .DOUT(N__21784),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__21786),
            .PADOUT(N__21785),
            .PADIN(N__21784),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__21777),
            .DIN(N__21776),
            .DOUT(N__21775),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__21777),
            .PADOUT(N__21776),
            .PADIN(N__21775),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21416),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__21768),
            .DIN(N__21767),
            .DOUT(N__21766),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__21768),
            .PADOUT(N__21767),
            .PADIN(N__21766),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__21759),
            .DIN(N__21758),
            .DOUT(N__21757),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__21759),
            .PADOUT(N__21758),
            .PADIN(N__21757),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__21750),
            .DIN(N__21749),
            .DOUT(N__21748),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__21750),
            .PADOUT(N__21749),
            .PADIN(N__21748),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__21741),
            .DIN(N__21740),
            .DOUT(N__21739),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__21741),
            .PADOUT(N__21740),
            .PADIN(N__21739),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18950),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__21732),
            .DIN(N__21731),
            .DOUT(N__21730),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__21732),
            .PADOUT(N__21731),
            .PADIN(N__21730),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13892),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__21723),
            .DIN(N__21722),
            .DOUT(N__21721),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__21723),
            .PADOUT(N__21722),
            .PADIN(N__21721),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__21714),
            .DIN(N__21713),
            .DOUT(N__21712),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__21714),
            .PADOUT(N__21713),
            .PADIN(N__21712),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15176),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__21705),
            .DIN(N__21704),
            .DOUT(N__21703),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__21705),
            .PADOUT(N__21704),
            .PADIN(N__21703),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5172 (
            .O(N__21686),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__5171 (
            .O(N__21683),
            .I(N__21672));
    InMux I__5170 (
            .O(N__21682),
            .I(N__21667));
    InMux I__5169 (
            .O(N__21681),
            .I(N__21661));
    InMux I__5168 (
            .O(N__21680),
            .I(N__21658));
    InMux I__5167 (
            .O(N__21679),
            .I(N__21653));
    InMux I__5166 (
            .O(N__21678),
            .I(N__21653));
    InMux I__5165 (
            .O(N__21677),
            .I(N__21646));
    InMux I__5164 (
            .O(N__21676),
            .I(N__21646));
    InMux I__5163 (
            .O(N__21675),
            .I(N__21646));
    InMux I__5162 (
            .O(N__21672),
            .I(N__21639));
    InMux I__5161 (
            .O(N__21671),
            .I(N__21639));
    InMux I__5160 (
            .O(N__21670),
            .I(N__21639));
    LocalMux I__5159 (
            .O(N__21667),
            .I(N__21636));
    InMux I__5158 (
            .O(N__21666),
            .I(N__21633));
    InMux I__5157 (
            .O(N__21665),
            .I(N__21628));
    InMux I__5156 (
            .O(N__21664),
            .I(N__21628));
    LocalMux I__5155 (
            .O(N__21661),
            .I(N__21625));
    LocalMux I__5154 (
            .O(N__21658),
            .I(N__21620));
    LocalMux I__5153 (
            .O(N__21653),
            .I(N__21620));
    LocalMux I__5152 (
            .O(N__21646),
            .I(N__21609));
    LocalMux I__5151 (
            .O(N__21639),
            .I(N__21609));
    Span4Mux_v I__5150 (
            .O(N__21636),
            .I(N__21609));
    LocalMux I__5149 (
            .O(N__21633),
            .I(N__21609));
    LocalMux I__5148 (
            .O(N__21628),
            .I(N__21609));
    Span4Mux_h I__5147 (
            .O(N__21625),
            .I(N__21606));
    Span4Mux_v I__5146 (
            .O(N__21620),
            .I(N__21601));
    Span4Mux_v I__5145 (
            .O(N__21609),
            .I(N__21601));
    Odrv4 I__5144 (
            .O(N__21606),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__5143 (
            .O(N__21601),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    CEMux I__5142 (
            .O(N__21596),
            .I(N__21581));
    CEMux I__5141 (
            .O(N__21595),
            .I(N__21581));
    CEMux I__5140 (
            .O(N__21594),
            .I(N__21581));
    CEMux I__5139 (
            .O(N__21593),
            .I(N__21581));
    CEMux I__5138 (
            .O(N__21592),
            .I(N__21581));
    GlobalMux I__5137 (
            .O(N__21581),
            .I(N__21578));
    gio2CtrlBuf I__5136 (
            .O(N__21578),
            .I(\delay_measurement_inst.delay_tr_timer.N_180_i_g ));
    InMux I__5135 (
            .O(N__21575),
            .I(N__21572));
    LocalMux I__5134 (
            .O(N__21572),
            .I(N__21568));
    InMux I__5133 (
            .O(N__21571),
            .I(N__21565));
    Span4Mux_s1_v I__5132 (
            .O(N__21568),
            .I(N__21560));
    LocalMux I__5131 (
            .O(N__21565),
            .I(N__21560));
    Span4Mux_v I__5130 (
            .O(N__21560),
            .I(N__21557));
    Span4Mux_h I__5129 (
            .O(N__21557),
            .I(N__21551));
    InMux I__5128 (
            .O(N__21556),
            .I(N__21548));
    CascadeMux I__5127 (
            .O(N__21555),
            .I(N__21545));
    InMux I__5126 (
            .O(N__21554),
            .I(N__21542));
    Span4Mux_v I__5125 (
            .O(N__21551),
            .I(N__21537));
    LocalMux I__5124 (
            .O(N__21548),
            .I(N__21537));
    InMux I__5123 (
            .O(N__21545),
            .I(N__21534));
    LocalMux I__5122 (
            .O(N__21542),
            .I(N__21531));
    Span4Mux_v I__5121 (
            .O(N__21537),
            .I(N__21527));
    LocalMux I__5120 (
            .O(N__21534),
            .I(N__21524));
    Span4Mux_v I__5119 (
            .O(N__21531),
            .I(N__21521));
    InMux I__5118 (
            .O(N__21530),
            .I(N__21518));
    Sp12to4 I__5117 (
            .O(N__21527),
            .I(N__21513));
    Span12Mux_s6_h I__5116 (
            .O(N__21524),
            .I(N__21513));
    Span4Mux_h I__5115 (
            .O(N__21521),
            .I(N__21510));
    LocalMux I__5114 (
            .O(N__21518),
            .I(N__21507));
    Span12Mux_v I__5113 (
            .O(N__21513),
            .I(N__21504));
    Sp12to4 I__5112 (
            .O(N__21510),
            .I(N__21499));
    Span12Mux_h I__5111 (
            .O(N__21507),
            .I(N__21499));
    Span12Mux_h I__5110 (
            .O(N__21504),
            .I(N__21496));
    Span12Mux_v I__5109 (
            .O(N__21499),
            .I(N__21493));
    Odrv12 I__5108 (
            .O(N__21496),
            .I(start_stop_c));
    Odrv12 I__5107 (
            .O(N__21493),
            .I(start_stop_c));
    CascadeMux I__5106 (
            .O(N__21488),
            .I(N__21484));
    InMux I__5105 (
            .O(N__21487),
            .I(N__21481));
    InMux I__5104 (
            .O(N__21484),
            .I(N__21477));
    LocalMux I__5103 (
            .O(N__21481),
            .I(N__21474));
    InMux I__5102 (
            .O(N__21480),
            .I(N__21471));
    LocalMux I__5101 (
            .O(N__21477),
            .I(N__21468));
    Span4Mux_v I__5100 (
            .O(N__21474),
            .I(N__21465));
    LocalMux I__5099 (
            .O(N__21471),
            .I(N__21460));
    Span4Mux_v I__5098 (
            .O(N__21468),
            .I(N__21455));
    Span4Mux_h I__5097 (
            .O(N__21465),
            .I(N__21455));
    InMux I__5096 (
            .O(N__21464),
            .I(N__21452));
    InMux I__5095 (
            .O(N__21463),
            .I(N__21449));
    Odrv12 I__5094 (
            .O(N__21460),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    Odrv4 I__5093 (
            .O(N__21455),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__5092 (
            .O(N__21452),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__5091 (
            .O(N__21449),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    InMux I__5090 (
            .O(N__21440),
            .I(N__21437));
    LocalMux I__5089 (
            .O(N__21437),
            .I(\phase_controller_inst1.N_110 ));
    InMux I__5088 (
            .O(N__21434),
            .I(N__21431));
    LocalMux I__5087 (
            .O(N__21431),
            .I(N__21428));
    Span4Mux_v I__5086 (
            .O(N__21428),
            .I(N__21425));
    Odrv4 I__5085 (
            .O(N__21425),
            .I(delay_tr_input_c));
    InMux I__5084 (
            .O(N__21422),
            .I(N__21419));
    LocalMux I__5083 (
            .O(N__21419),
            .I(delay_tr_d1));
    IoInMux I__5082 (
            .O(N__21416),
            .I(N__21413));
    LocalMux I__5081 (
            .O(N__21413),
            .I(N__21410));
    Span4Mux_s3_v I__5080 (
            .O(N__21410),
            .I(N__21407));
    Span4Mux_h I__5079 (
            .O(N__21407),
            .I(N__21404));
    Sp12to4 I__5078 (
            .O(N__21404),
            .I(N__21401));
    Span12Mux_v I__5077 (
            .O(N__21401),
            .I(N__21397));
    InMux I__5076 (
            .O(N__21400),
            .I(N__21394));
    Odrv12 I__5075 (
            .O(N__21397),
            .I(T23_c));
    LocalMux I__5074 (
            .O(N__21394),
            .I(T23_c));
    CascadeMux I__5073 (
            .O(N__21389),
            .I(N__21384));
    CascadeMux I__5072 (
            .O(N__21388),
            .I(N__21381));
    CascadeMux I__5071 (
            .O(N__21387),
            .I(N__21378));
    InMux I__5070 (
            .O(N__21384),
            .I(N__21360));
    InMux I__5069 (
            .O(N__21381),
            .I(N__21360));
    InMux I__5068 (
            .O(N__21378),
            .I(N__21360));
    InMux I__5067 (
            .O(N__21377),
            .I(N__21357));
    InMux I__5066 (
            .O(N__21376),
            .I(N__21354));
    InMux I__5065 (
            .O(N__21375),
            .I(N__21351));
    CascadeMux I__5064 (
            .O(N__21374),
            .I(N__21340));
    InMux I__5063 (
            .O(N__21373),
            .I(N__21323));
    InMux I__5062 (
            .O(N__21372),
            .I(N__21323));
    InMux I__5061 (
            .O(N__21371),
            .I(N__21323));
    InMux I__5060 (
            .O(N__21370),
            .I(N__21323));
    InMux I__5059 (
            .O(N__21369),
            .I(N__21323));
    InMux I__5058 (
            .O(N__21368),
            .I(N__21323));
    InMux I__5057 (
            .O(N__21367),
            .I(N__21323));
    LocalMux I__5056 (
            .O(N__21360),
            .I(N__21318));
    LocalMux I__5055 (
            .O(N__21357),
            .I(N__21318));
    LocalMux I__5054 (
            .O(N__21354),
            .I(N__21313));
    LocalMux I__5053 (
            .O(N__21351),
            .I(N__21313));
    InMux I__5052 (
            .O(N__21350),
            .I(N__21300));
    InMux I__5051 (
            .O(N__21349),
            .I(N__21300));
    InMux I__5050 (
            .O(N__21348),
            .I(N__21300));
    InMux I__5049 (
            .O(N__21347),
            .I(N__21300));
    InMux I__5048 (
            .O(N__21346),
            .I(N__21300));
    InMux I__5047 (
            .O(N__21345),
            .I(N__21287));
    InMux I__5046 (
            .O(N__21344),
            .I(N__21287));
    InMux I__5045 (
            .O(N__21343),
            .I(N__21287));
    InMux I__5044 (
            .O(N__21340),
            .I(N__21287));
    InMux I__5043 (
            .O(N__21339),
            .I(N__21287));
    InMux I__5042 (
            .O(N__21338),
            .I(N__21287));
    LocalMux I__5041 (
            .O(N__21323),
            .I(N__21282));
    Span4Mux_h I__5040 (
            .O(N__21318),
            .I(N__21282));
    Span4Mux_v I__5039 (
            .O(N__21313),
            .I(N__21279));
    InMux I__5038 (
            .O(N__21312),
            .I(N__21274));
    InMux I__5037 (
            .O(N__21311),
            .I(N__21274));
    LocalMux I__5036 (
            .O(N__21300),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__5035 (
            .O(N__21287),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__5034 (
            .O(N__21282),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__5033 (
            .O(N__21279),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__5032 (
            .O(N__21274),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__5031 (
            .O(N__21263),
            .I(N__21260));
    InMux I__5030 (
            .O(N__21260),
            .I(N__21257));
    LocalMux I__5029 (
            .O(N__21257),
            .I(\phase_controller_inst1.stoper_hc.N_60 ));
    InMux I__5028 (
            .O(N__21254),
            .I(N__21251));
    LocalMux I__5027 (
            .O(N__21251),
            .I(N__21243));
    InMux I__5026 (
            .O(N__21250),
            .I(N__21232));
    InMux I__5025 (
            .O(N__21249),
            .I(N__21232));
    InMux I__5024 (
            .O(N__21248),
            .I(N__21232));
    InMux I__5023 (
            .O(N__21247),
            .I(N__21232));
    InMux I__5022 (
            .O(N__21246),
            .I(N__21232));
    Odrv12 I__5021 (
            .O(N__21243),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__5020 (
            .O(N__21232),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__5019 (
            .O(N__21227),
            .I(N__21223));
    InMux I__5018 (
            .O(N__21226),
            .I(N__21220));
    LocalMux I__5017 (
            .O(N__21223),
            .I(N__21215));
    LocalMux I__5016 (
            .O(N__21220),
            .I(N__21215));
    Span4Mux_h I__5015 (
            .O(N__21215),
            .I(N__21211));
    InMux I__5014 (
            .O(N__21214),
            .I(N__21207));
    Span4Mux_v I__5013 (
            .O(N__21211),
            .I(N__21204));
    InMux I__5012 (
            .O(N__21210),
            .I(N__21201));
    LocalMux I__5011 (
            .O(N__21207),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__5010 (
            .O(N__21204),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5009 (
            .O(N__21201),
            .I(\phase_controller_inst1.hc_time_passed ));
    ClkMux I__5008 (
            .O(N__21194),
            .I(N__20906));
    ClkMux I__5007 (
            .O(N__21193),
            .I(N__20906));
    ClkMux I__5006 (
            .O(N__21192),
            .I(N__20906));
    ClkMux I__5005 (
            .O(N__21191),
            .I(N__20906));
    ClkMux I__5004 (
            .O(N__21190),
            .I(N__20906));
    ClkMux I__5003 (
            .O(N__21189),
            .I(N__20906));
    ClkMux I__5002 (
            .O(N__21188),
            .I(N__20906));
    ClkMux I__5001 (
            .O(N__21187),
            .I(N__20906));
    ClkMux I__5000 (
            .O(N__21186),
            .I(N__20906));
    ClkMux I__4999 (
            .O(N__21185),
            .I(N__20906));
    ClkMux I__4998 (
            .O(N__21184),
            .I(N__20906));
    ClkMux I__4997 (
            .O(N__21183),
            .I(N__20906));
    ClkMux I__4996 (
            .O(N__21182),
            .I(N__20906));
    ClkMux I__4995 (
            .O(N__21181),
            .I(N__20906));
    ClkMux I__4994 (
            .O(N__21180),
            .I(N__20906));
    ClkMux I__4993 (
            .O(N__21179),
            .I(N__20906));
    ClkMux I__4992 (
            .O(N__21178),
            .I(N__20906));
    ClkMux I__4991 (
            .O(N__21177),
            .I(N__20906));
    ClkMux I__4990 (
            .O(N__21176),
            .I(N__20906));
    ClkMux I__4989 (
            .O(N__21175),
            .I(N__20906));
    ClkMux I__4988 (
            .O(N__21174),
            .I(N__20906));
    ClkMux I__4987 (
            .O(N__21173),
            .I(N__20906));
    ClkMux I__4986 (
            .O(N__21172),
            .I(N__20906));
    ClkMux I__4985 (
            .O(N__21171),
            .I(N__20906));
    ClkMux I__4984 (
            .O(N__21170),
            .I(N__20906));
    ClkMux I__4983 (
            .O(N__21169),
            .I(N__20906));
    ClkMux I__4982 (
            .O(N__21168),
            .I(N__20906));
    ClkMux I__4981 (
            .O(N__21167),
            .I(N__20906));
    ClkMux I__4980 (
            .O(N__21166),
            .I(N__20906));
    ClkMux I__4979 (
            .O(N__21165),
            .I(N__20906));
    ClkMux I__4978 (
            .O(N__21164),
            .I(N__20906));
    ClkMux I__4977 (
            .O(N__21163),
            .I(N__20906));
    ClkMux I__4976 (
            .O(N__21162),
            .I(N__20906));
    ClkMux I__4975 (
            .O(N__21161),
            .I(N__20906));
    ClkMux I__4974 (
            .O(N__21160),
            .I(N__20906));
    ClkMux I__4973 (
            .O(N__21159),
            .I(N__20906));
    ClkMux I__4972 (
            .O(N__21158),
            .I(N__20906));
    ClkMux I__4971 (
            .O(N__21157),
            .I(N__20906));
    ClkMux I__4970 (
            .O(N__21156),
            .I(N__20906));
    ClkMux I__4969 (
            .O(N__21155),
            .I(N__20906));
    ClkMux I__4968 (
            .O(N__21154),
            .I(N__20906));
    ClkMux I__4967 (
            .O(N__21153),
            .I(N__20906));
    ClkMux I__4966 (
            .O(N__21152),
            .I(N__20906));
    ClkMux I__4965 (
            .O(N__21151),
            .I(N__20906));
    ClkMux I__4964 (
            .O(N__21150),
            .I(N__20906));
    ClkMux I__4963 (
            .O(N__21149),
            .I(N__20906));
    ClkMux I__4962 (
            .O(N__21148),
            .I(N__20906));
    ClkMux I__4961 (
            .O(N__21147),
            .I(N__20906));
    ClkMux I__4960 (
            .O(N__21146),
            .I(N__20906));
    ClkMux I__4959 (
            .O(N__21145),
            .I(N__20906));
    ClkMux I__4958 (
            .O(N__21144),
            .I(N__20906));
    ClkMux I__4957 (
            .O(N__21143),
            .I(N__20906));
    ClkMux I__4956 (
            .O(N__21142),
            .I(N__20906));
    ClkMux I__4955 (
            .O(N__21141),
            .I(N__20906));
    ClkMux I__4954 (
            .O(N__21140),
            .I(N__20906));
    ClkMux I__4953 (
            .O(N__21139),
            .I(N__20906));
    ClkMux I__4952 (
            .O(N__21138),
            .I(N__20906));
    ClkMux I__4951 (
            .O(N__21137),
            .I(N__20906));
    ClkMux I__4950 (
            .O(N__21136),
            .I(N__20906));
    ClkMux I__4949 (
            .O(N__21135),
            .I(N__20906));
    ClkMux I__4948 (
            .O(N__21134),
            .I(N__20906));
    ClkMux I__4947 (
            .O(N__21133),
            .I(N__20906));
    ClkMux I__4946 (
            .O(N__21132),
            .I(N__20906));
    ClkMux I__4945 (
            .O(N__21131),
            .I(N__20906));
    ClkMux I__4944 (
            .O(N__21130),
            .I(N__20906));
    ClkMux I__4943 (
            .O(N__21129),
            .I(N__20906));
    ClkMux I__4942 (
            .O(N__21128),
            .I(N__20906));
    ClkMux I__4941 (
            .O(N__21127),
            .I(N__20906));
    ClkMux I__4940 (
            .O(N__21126),
            .I(N__20906));
    ClkMux I__4939 (
            .O(N__21125),
            .I(N__20906));
    ClkMux I__4938 (
            .O(N__21124),
            .I(N__20906));
    ClkMux I__4937 (
            .O(N__21123),
            .I(N__20906));
    ClkMux I__4936 (
            .O(N__21122),
            .I(N__20906));
    ClkMux I__4935 (
            .O(N__21121),
            .I(N__20906));
    ClkMux I__4934 (
            .O(N__21120),
            .I(N__20906));
    ClkMux I__4933 (
            .O(N__21119),
            .I(N__20906));
    ClkMux I__4932 (
            .O(N__21118),
            .I(N__20906));
    ClkMux I__4931 (
            .O(N__21117),
            .I(N__20906));
    ClkMux I__4930 (
            .O(N__21116),
            .I(N__20906));
    ClkMux I__4929 (
            .O(N__21115),
            .I(N__20906));
    ClkMux I__4928 (
            .O(N__21114),
            .I(N__20906));
    ClkMux I__4927 (
            .O(N__21113),
            .I(N__20906));
    ClkMux I__4926 (
            .O(N__21112),
            .I(N__20906));
    ClkMux I__4925 (
            .O(N__21111),
            .I(N__20906));
    ClkMux I__4924 (
            .O(N__21110),
            .I(N__20906));
    ClkMux I__4923 (
            .O(N__21109),
            .I(N__20906));
    ClkMux I__4922 (
            .O(N__21108),
            .I(N__20906));
    ClkMux I__4921 (
            .O(N__21107),
            .I(N__20906));
    ClkMux I__4920 (
            .O(N__21106),
            .I(N__20906));
    ClkMux I__4919 (
            .O(N__21105),
            .I(N__20906));
    ClkMux I__4918 (
            .O(N__21104),
            .I(N__20906));
    ClkMux I__4917 (
            .O(N__21103),
            .I(N__20906));
    ClkMux I__4916 (
            .O(N__21102),
            .I(N__20906));
    ClkMux I__4915 (
            .O(N__21101),
            .I(N__20906));
    ClkMux I__4914 (
            .O(N__21100),
            .I(N__20906));
    ClkMux I__4913 (
            .O(N__21099),
            .I(N__20906));
    GlobalMux I__4912 (
            .O(N__20906),
            .I(clk_100mhz));
    CascadeMux I__4911 (
            .O(N__20903),
            .I(N__20895));
    InMux I__4910 (
            .O(N__20902),
            .I(N__20886));
    InMux I__4909 (
            .O(N__20901),
            .I(N__20883));
    InMux I__4908 (
            .O(N__20900),
            .I(N__20880));
    InMux I__4907 (
            .O(N__20899),
            .I(N__20877));
    InMux I__4906 (
            .O(N__20898),
            .I(N__20874));
    InMux I__4905 (
            .O(N__20895),
            .I(N__20869));
    InMux I__4904 (
            .O(N__20894),
            .I(N__20869));
    InMux I__4903 (
            .O(N__20893),
            .I(N__20866));
    InMux I__4902 (
            .O(N__20892),
            .I(N__20863));
    InMux I__4901 (
            .O(N__20891),
            .I(N__20856));
    InMux I__4900 (
            .O(N__20890),
            .I(N__20856));
    InMux I__4899 (
            .O(N__20889),
            .I(N__20856));
    LocalMux I__4898 (
            .O(N__20886),
            .I(N__20853));
    LocalMux I__4897 (
            .O(N__20883),
            .I(N__20850));
    LocalMux I__4896 (
            .O(N__20880),
            .I(N__20847));
    LocalMux I__4895 (
            .O(N__20877),
            .I(N__20840));
    LocalMux I__4894 (
            .O(N__20874),
            .I(N__20815));
    LocalMux I__4893 (
            .O(N__20869),
            .I(N__20773));
    LocalMux I__4892 (
            .O(N__20866),
            .I(N__20770));
    LocalMux I__4891 (
            .O(N__20863),
            .I(N__20766));
    LocalMux I__4890 (
            .O(N__20856),
            .I(N__20763));
    Glb2LocalMux I__4889 (
            .O(N__20853),
            .I(N__20597));
    Glb2LocalMux I__4888 (
            .O(N__20850),
            .I(N__20597));
    Glb2LocalMux I__4887 (
            .O(N__20847),
            .I(N__20597));
    SRMux I__4886 (
            .O(N__20846),
            .I(N__20597));
    SRMux I__4885 (
            .O(N__20845),
            .I(N__20597));
    SRMux I__4884 (
            .O(N__20844),
            .I(N__20597));
    SRMux I__4883 (
            .O(N__20843),
            .I(N__20597));
    Glb2LocalMux I__4882 (
            .O(N__20840),
            .I(N__20597));
    SRMux I__4881 (
            .O(N__20839),
            .I(N__20597));
    SRMux I__4880 (
            .O(N__20838),
            .I(N__20597));
    SRMux I__4879 (
            .O(N__20837),
            .I(N__20597));
    SRMux I__4878 (
            .O(N__20836),
            .I(N__20597));
    SRMux I__4877 (
            .O(N__20835),
            .I(N__20597));
    SRMux I__4876 (
            .O(N__20834),
            .I(N__20597));
    SRMux I__4875 (
            .O(N__20833),
            .I(N__20597));
    SRMux I__4874 (
            .O(N__20832),
            .I(N__20597));
    SRMux I__4873 (
            .O(N__20831),
            .I(N__20597));
    SRMux I__4872 (
            .O(N__20830),
            .I(N__20597));
    SRMux I__4871 (
            .O(N__20829),
            .I(N__20597));
    SRMux I__4870 (
            .O(N__20828),
            .I(N__20597));
    SRMux I__4869 (
            .O(N__20827),
            .I(N__20597));
    SRMux I__4868 (
            .O(N__20826),
            .I(N__20597));
    SRMux I__4867 (
            .O(N__20825),
            .I(N__20597));
    SRMux I__4866 (
            .O(N__20824),
            .I(N__20597));
    SRMux I__4865 (
            .O(N__20823),
            .I(N__20597));
    SRMux I__4864 (
            .O(N__20822),
            .I(N__20597));
    SRMux I__4863 (
            .O(N__20821),
            .I(N__20597));
    SRMux I__4862 (
            .O(N__20820),
            .I(N__20597));
    SRMux I__4861 (
            .O(N__20819),
            .I(N__20597));
    SRMux I__4860 (
            .O(N__20818),
            .I(N__20597));
    Glb2LocalMux I__4859 (
            .O(N__20815),
            .I(N__20597));
    SRMux I__4858 (
            .O(N__20814),
            .I(N__20597));
    SRMux I__4857 (
            .O(N__20813),
            .I(N__20597));
    SRMux I__4856 (
            .O(N__20812),
            .I(N__20597));
    SRMux I__4855 (
            .O(N__20811),
            .I(N__20597));
    SRMux I__4854 (
            .O(N__20810),
            .I(N__20597));
    SRMux I__4853 (
            .O(N__20809),
            .I(N__20597));
    SRMux I__4852 (
            .O(N__20808),
            .I(N__20597));
    SRMux I__4851 (
            .O(N__20807),
            .I(N__20597));
    SRMux I__4850 (
            .O(N__20806),
            .I(N__20597));
    SRMux I__4849 (
            .O(N__20805),
            .I(N__20597));
    SRMux I__4848 (
            .O(N__20804),
            .I(N__20597));
    SRMux I__4847 (
            .O(N__20803),
            .I(N__20597));
    SRMux I__4846 (
            .O(N__20802),
            .I(N__20597));
    SRMux I__4845 (
            .O(N__20801),
            .I(N__20597));
    SRMux I__4844 (
            .O(N__20800),
            .I(N__20597));
    SRMux I__4843 (
            .O(N__20799),
            .I(N__20597));
    SRMux I__4842 (
            .O(N__20798),
            .I(N__20597));
    SRMux I__4841 (
            .O(N__20797),
            .I(N__20597));
    SRMux I__4840 (
            .O(N__20796),
            .I(N__20597));
    SRMux I__4839 (
            .O(N__20795),
            .I(N__20597));
    SRMux I__4838 (
            .O(N__20794),
            .I(N__20597));
    SRMux I__4837 (
            .O(N__20793),
            .I(N__20597));
    SRMux I__4836 (
            .O(N__20792),
            .I(N__20597));
    SRMux I__4835 (
            .O(N__20791),
            .I(N__20597));
    SRMux I__4834 (
            .O(N__20790),
            .I(N__20597));
    SRMux I__4833 (
            .O(N__20789),
            .I(N__20597));
    SRMux I__4832 (
            .O(N__20788),
            .I(N__20597));
    SRMux I__4831 (
            .O(N__20787),
            .I(N__20597));
    SRMux I__4830 (
            .O(N__20786),
            .I(N__20597));
    SRMux I__4829 (
            .O(N__20785),
            .I(N__20597));
    SRMux I__4828 (
            .O(N__20784),
            .I(N__20597));
    SRMux I__4827 (
            .O(N__20783),
            .I(N__20597));
    SRMux I__4826 (
            .O(N__20782),
            .I(N__20597));
    SRMux I__4825 (
            .O(N__20781),
            .I(N__20597));
    SRMux I__4824 (
            .O(N__20780),
            .I(N__20597));
    SRMux I__4823 (
            .O(N__20779),
            .I(N__20597));
    SRMux I__4822 (
            .O(N__20778),
            .I(N__20597));
    SRMux I__4821 (
            .O(N__20777),
            .I(N__20597));
    SRMux I__4820 (
            .O(N__20776),
            .I(N__20597));
    Glb2LocalMux I__4819 (
            .O(N__20773),
            .I(N__20597));
    Glb2LocalMux I__4818 (
            .O(N__20770),
            .I(N__20597));
    SRMux I__4817 (
            .O(N__20769),
            .I(N__20597));
    Glb2LocalMux I__4816 (
            .O(N__20766),
            .I(N__20597));
    Glb2LocalMux I__4815 (
            .O(N__20763),
            .I(N__20597));
    SRMux I__4814 (
            .O(N__20762),
            .I(N__20597));
    SRMux I__4813 (
            .O(N__20761),
            .I(N__20597));
    SRMux I__4812 (
            .O(N__20760),
            .I(N__20597));
    SRMux I__4811 (
            .O(N__20759),
            .I(N__20597));
    SRMux I__4810 (
            .O(N__20758),
            .I(N__20597));
    GlobalMux I__4809 (
            .O(N__20597),
            .I(N__20594));
    gio2CtrlBuf I__4808 (
            .O(N__20594),
            .I(red_c_g));
    CascadeMux I__4807 (
            .O(N__20591),
            .I(N__20586));
    InMux I__4806 (
            .O(N__20590),
            .I(N__20583));
    InMux I__4805 (
            .O(N__20589),
            .I(N__20580));
    InMux I__4804 (
            .O(N__20586),
            .I(N__20577));
    LocalMux I__4803 (
            .O(N__20583),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__4802 (
            .O(N__20580),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__4801 (
            .O(N__20577),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    CascadeMux I__4800 (
            .O(N__20570),
            .I(N__20567));
    InMux I__4799 (
            .O(N__20567),
            .I(N__20564));
    LocalMux I__4798 (
            .O(N__20564),
            .I(N__20561));
    Odrv4 I__4797 (
            .O(N__20561),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__4796 (
            .O(N__20558),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__4795 (
            .O(N__20555),
            .I(N__20550));
    InMux I__4794 (
            .O(N__20554),
            .I(N__20547));
    InMux I__4793 (
            .O(N__20553),
            .I(N__20544));
    InMux I__4792 (
            .O(N__20550),
            .I(N__20541));
    LocalMux I__4791 (
            .O(N__20547),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__4790 (
            .O(N__20544),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__4789 (
            .O(N__20541),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__4788 (
            .O(N__20534),
            .I(N__20531));
    LocalMux I__4787 (
            .O(N__20531),
            .I(N__20528));
    Span4Mux_h I__4786 (
            .O(N__20528),
            .I(N__20525));
    Odrv4 I__4785 (
            .O(N__20525),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__4784 (
            .O(N__20522),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__4783 (
            .O(N__20519),
            .I(N__20514));
    InMux I__4782 (
            .O(N__20518),
            .I(N__20511));
    InMux I__4781 (
            .O(N__20517),
            .I(N__20508));
    InMux I__4780 (
            .O(N__20514),
            .I(N__20505));
    LocalMux I__4779 (
            .O(N__20511),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__4778 (
            .O(N__20508),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__4777 (
            .O(N__20505),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__4776 (
            .O(N__20498),
            .I(N__20495));
    LocalMux I__4775 (
            .O(N__20495),
            .I(N__20492));
    Odrv4 I__4774 (
            .O(N__20492),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__4773 (
            .O(N__20489),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__4772 (
            .O(N__20486),
            .I(N__20481));
    InMux I__4771 (
            .O(N__20485),
            .I(N__20478));
    InMux I__4770 (
            .O(N__20484),
            .I(N__20475));
    InMux I__4769 (
            .O(N__20481),
            .I(N__20472));
    LocalMux I__4768 (
            .O(N__20478),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__4767 (
            .O(N__20475),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__4766 (
            .O(N__20472),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__4765 (
            .O(N__20465),
            .I(N__20462));
    LocalMux I__4764 (
            .O(N__20462),
            .I(N__20459));
    Odrv4 I__4763 (
            .O(N__20459),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__4762 (
            .O(N__20456),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__4761 (
            .O(N__20453),
            .I(N__20448));
    InMux I__4760 (
            .O(N__20452),
            .I(N__20445));
    InMux I__4759 (
            .O(N__20451),
            .I(N__20442));
    InMux I__4758 (
            .O(N__20448),
            .I(N__20439));
    LocalMux I__4757 (
            .O(N__20445),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__4756 (
            .O(N__20442),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__4755 (
            .O(N__20439),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__4754 (
            .O(N__20432),
            .I(N__20429));
    LocalMux I__4753 (
            .O(N__20429),
            .I(N__20426));
    Span4Mux_v I__4752 (
            .O(N__20426),
            .I(N__20423));
    Odrv4 I__4751 (
            .O(N__20423),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__4750 (
            .O(N__20420),
            .I(bfn_13_22_0_));
    CascadeMux I__4749 (
            .O(N__20417),
            .I(N__20412));
    InMux I__4748 (
            .O(N__20416),
            .I(N__20409));
    InMux I__4747 (
            .O(N__20415),
            .I(N__20406));
    InMux I__4746 (
            .O(N__20412),
            .I(N__20403));
    LocalMux I__4745 (
            .O(N__20409),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__4744 (
            .O(N__20406),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__4743 (
            .O(N__20403),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    CascadeMux I__4742 (
            .O(N__20396),
            .I(N__20393));
    InMux I__4741 (
            .O(N__20393),
            .I(N__20390));
    LocalMux I__4740 (
            .O(N__20390),
            .I(N__20387));
    Span4Mux_v I__4739 (
            .O(N__20387),
            .I(N__20384));
    Odrv4 I__4738 (
            .O(N__20384),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__4737 (
            .O(N__20381),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    CascadeMux I__4736 (
            .O(N__20378),
            .I(N__20373));
    InMux I__4735 (
            .O(N__20377),
            .I(N__20370));
    InMux I__4734 (
            .O(N__20376),
            .I(N__20367));
    InMux I__4733 (
            .O(N__20373),
            .I(N__20364));
    LocalMux I__4732 (
            .O(N__20370),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__4731 (
            .O(N__20367),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__4730 (
            .O(N__20364),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    CascadeMux I__4729 (
            .O(N__20357),
            .I(N__20353));
    InMux I__4728 (
            .O(N__20356),
            .I(N__20350));
    InMux I__4727 (
            .O(N__20353),
            .I(N__20347));
    LocalMux I__4726 (
            .O(N__20350),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__4725 (
            .O(N__20347),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__4724 (
            .O(N__20342),
            .I(N__20339));
    LocalMux I__4723 (
            .O(N__20339),
            .I(N__20336));
    Odrv4 I__4722 (
            .O(N__20336),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__4721 (
            .O(N__20333),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__4720 (
            .O(N__20330),
            .I(N__20325));
    InMux I__4719 (
            .O(N__20329),
            .I(N__20322));
    InMux I__4718 (
            .O(N__20328),
            .I(N__20319));
    InMux I__4717 (
            .O(N__20325),
            .I(N__20316));
    LocalMux I__4716 (
            .O(N__20322),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__4715 (
            .O(N__20319),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__4714 (
            .O(N__20316),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    CascadeMux I__4713 (
            .O(N__20309),
            .I(N__20305));
    InMux I__4712 (
            .O(N__20308),
            .I(N__20302));
    InMux I__4711 (
            .O(N__20305),
            .I(N__20299));
    LocalMux I__4710 (
            .O(N__20302),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__4709 (
            .O(N__20299),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    InMux I__4708 (
            .O(N__20294),
            .I(N__20291));
    LocalMux I__4707 (
            .O(N__20291),
            .I(N__20288));
    Odrv4 I__4706 (
            .O(N__20288),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__4705 (
            .O(N__20285),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    CascadeMux I__4704 (
            .O(N__20282),
            .I(N__20277));
    InMux I__4703 (
            .O(N__20281),
            .I(N__20274));
    InMux I__4702 (
            .O(N__20280),
            .I(N__20271));
    InMux I__4701 (
            .O(N__20277),
            .I(N__20268));
    LocalMux I__4700 (
            .O(N__20274),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__4699 (
            .O(N__20271),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__4698 (
            .O(N__20268),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    CascadeMux I__4697 (
            .O(N__20261),
            .I(N__20253));
    InMux I__4696 (
            .O(N__20260),
            .I(N__20250));
    InMux I__4695 (
            .O(N__20259),
            .I(N__20247));
    InMux I__4694 (
            .O(N__20258),
            .I(N__20240));
    InMux I__4693 (
            .O(N__20257),
            .I(N__20240));
    InMux I__4692 (
            .O(N__20256),
            .I(N__20240));
    InMux I__4691 (
            .O(N__20253),
            .I(N__20237));
    LocalMux I__4690 (
            .O(N__20250),
            .I(N__20232));
    LocalMux I__4689 (
            .O(N__20247),
            .I(N__20232));
    LocalMux I__4688 (
            .O(N__20240),
            .I(N__20229));
    LocalMux I__4687 (
            .O(N__20237),
            .I(N__20224));
    Span4Mux_v I__4686 (
            .O(N__20232),
            .I(N__20224));
    Span4Mux_v I__4685 (
            .O(N__20229),
            .I(N__20221));
    Span4Mux_h I__4684 (
            .O(N__20224),
            .I(N__20218));
    Odrv4 I__4683 (
            .O(N__20221),
            .I(\delay_measurement_inst.elapsed_time_tr_15 ));
    Odrv4 I__4682 (
            .O(N__20218),
            .I(\delay_measurement_inst.elapsed_time_tr_15 ));
    InMux I__4681 (
            .O(N__20213),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__4680 (
            .O(N__20210),
            .I(N__20205));
    InMux I__4679 (
            .O(N__20209),
            .I(N__20202));
    InMux I__4678 (
            .O(N__20208),
            .I(N__20199));
    InMux I__4677 (
            .O(N__20205),
            .I(N__20196));
    LocalMux I__4676 (
            .O(N__20202),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__4675 (
            .O(N__20199),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__4674 (
            .O(N__20196),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__4673 (
            .O(N__20189),
            .I(N__20184));
    InMux I__4672 (
            .O(N__20188),
            .I(N__20181));
    InMux I__4671 (
            .O(N__20187),
            .I(N__20178));
    LocalMux I__4670 (
            .O(N__20184),
            .I(N__20173));
    LocalMux I__4669 (
            .O(N__20181),
            .I(N__20173));
    LocalMux I__4668 (
            .O(N__20178),
            .I(N__20170));
    Span4Mux_v I__4667 (
            .O(N__20173),
            .I(N__20167));
    Span4Mux_v I__4666 (
            .O(N__20170),
            .I(N__20164));
    Span4Mux_h I__4665 (
            .O(N__20167),
            .I(N__20161));
    Odrv4 I__4664 (
            .O(N__20164),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    Odrv4 I__4663 (
            .O(N__20161),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__4662 (
            .O(N__20156),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__4661 (
            .O(N__20153),
            .I(N__20148));
    InMux I__4660 (
            .O(N__20152),
            .I(N__20145));
    InMux I__4659 (
            .O(N__20151),
            .I(N__20142));
    InMux I__4658 (
            .O(N__20148),
            .I(N__20139));
    LocalMux I__4657 (
            .O(N__20145),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__4656 (
            .O(N__20142),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__4655 (
            .O(N__20139),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__4654 (
            .O(N__20132),
            .I(N__20125));
    InMux I__4653 (
            .O(N__20131),
            .I(N__20125));
    InMux I__4652 (
            .O(N__20130),
            .I(N__20122));
    LocalMux I__4651 (
            .O(N__20125),
            .I(N__20119));
    LocalMux I__4650 (
            .O(N__20122),
            .I(N__20116));
    Span4Mux_h I__4649 (
            .O(N__20119),
            .I(N__20113));
    Odrv12 I__4648 (
            .O(N__20116),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv4 I__4647 (
            .O(N__20113),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__4646 (
            .O(N__20108),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__4645 (
            .O(N__20105),
            .I(N__20100));
    InMux I__4644 (
            .O(N__20104),
            .I(N__20097));
    InMux I__4643 (
            .O(N__20103),
            .I(N__20094));
    InMux I__4642 (
            .O(N__20100),
            .I(N__20091));
    LocalMux I__4641 (
            .O(N__20097),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__4640 (
            .O(N__20094),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__4639 (
            .O(N__20091),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    CascadeMux I__4638 (
            .O(N__20084),
            .I(N__20080));
    CascadeMux I__4637 (
            .O(N__20083),
            .I(N__20077));
    InMux I__4636 (
            .O(N__20080),
            .I(N__20073));
    InMux I__4635 (
            .O(N__20077),
            .I(N__20070));
    InMux I__4634 (
            .O(N__20076),
            .I(N__20067));
    LocalMux I__4633 (
            .O(N__20073),
            .I(N__20062));
    LocalMux I__4632 (
            .O(N__20070),
            .I(N__20062));
    LocalMux I__4631 (
            .O(N__20067),
            .I(N__20059));
    Span4Mux_h I__4630 (
            .O(N__20062),
            .I(N__20056));
    Odrv4 I__4629 (
            .O(N__20059),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv4 I__4628 (
            .O(N__20056),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    InMux I__4627 (
            .O(N__20051),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__4626 (
            .O(N__20048),
            .I(N__20043));
    InMux I__4625 (
            .O(N__20047),
            .I(N__20040));
    InMux I__4624 (
            .O(N__20046),
            .I(N__20037));
    InMux I__4623 (
            .O(N__20043),
            .I(N__20034));
    LocalMux I__4622 (
            .O(N__20040),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__4621 (
            .O(N__20037),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__4620 (
            .O(N__20034),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__4619 (
            .O(N__20027),
            .I(N__20023));
    CascadeMux I__4618 (
            .O(N__20026),
            .I(N__20019));
    LocalMux I__4617 (
            .O(N__20023),
            .I(N__20016));
    InMux I__4616 (
            .O(N__20022),
            .I(N__20011));
    InMux I__4615 (
            .O(N__20019),
            .I(N__20011));
    Span4Mux_v I__4614 (
            .O(N__20016),
            .I(N__20006));
    LocalMux I__4613 (
            .O(N__20011),
            .I(N__20006));
    Odrv4 I__4612 (
            .O(N__20006),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    InMux I__4611 (
            .O(N__20003),
            .I(bfn_13_21_0_));
    CascadeMux I__4610 (
            .O(N__20000),
            .I(N__19995));
    InMux I__4609 (
            .O(N__19999),
            .I(N__19992));
    InMux I__4608 (
            .O(N__19998),
            .I(N__19989));
    InMux I__4607 (
            .O(N__19995),
            .I(N__19986));
    LocalMux I__4606 (
            .O(N__19992),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__4605 (
            .O(N__19989),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__4604 (
            .O(N__19986),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    CascadeMux I__4603 (
            .O(N__19979),
            .I(N__19976));
    InMux I__4602 (
            .O(N__19976),
            .I(N__19973));
    LocalMux I__4601 (
            .O(N__19973),
            .I(N__19970));
    Odrv12 I__4600 (
            .O(N__19970),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__4599 (
            .O(N__19967),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__4598 (
            .O(N__19964),
            .I(N__19959));
    InMux I__4597 (
            .O(N__19963),
            .I(N__19956));
    InMux I__4596 (
            .O(N__19962),
            .I(N__19953));
    InMux I__4595 (
            .O(N__19959),
            .I(N__19950));
    LocalMux I__4594 (
            .O(N__19956),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__4593 (
            .O(N__19953),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__4592 (
            .O(N__19950),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__4591 (
            .O(N__19943),
            .I(N__19940));
    LocalMux I__4590 (
            .O(N__19940),
            .I(N__19937));
    Odrv4 I__4589 (
            .O(N__19937),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__4588 (
            .O(N__19934),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__4587 (
            .O(N__19931),
            .I(N__19926));
    InMux I__4586 (
            .O(N__19930),
            .I(N__19923));
    InMux I__4585 (
            .O(N__19929),
            .I(N__19920));
    InMux I__4584 (
            .O(N__19926),
            .I(N__19917));
    LocalMux I__4583 (
            .O(N__19923),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__4582 (
            .O(N__19920),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__4581 (
            .O(N__19917),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__4580 (
            .O(N__19910),
            .I(N__19907));
    LocalMux I__4579 (
            .O(N__19907),
            .I(N__19904));
    Odrv12 I__4578 (
            .O(N__19904),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__4577 (
            .O(N__19901),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__4576 (
            .O(N__19898),
            .I(N__19895));
    InMux I__4575 (
            .O(N__19895),
            .I(N__19892));
    LocalMux I__4574 (
            .O(N__19892),
            .I(N__19888));
    InMux I__4573 (
            .O(N__19891),
            .I(N__19885));
    Span4Mux_h I__4572 (
            .O(N__19888),
            .I(N__19882));
    LocalMux I__4571 (
            .O(N__19885),
            .I(N__19879));
    Odrv4 I__4570 (
            .O(N__19882),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    Odrv12 I__4569 (
            .O(N__19879),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__4568 (
            .O(N__19874),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__4567 (
            .O(N__19871),
            .I(N__19866));
    InMux I__4566 (
            .O(N__19870),
            .I(N__19863));
    InMux I__4565 (
            .O(N__19869),
            .I(N__19860));
    InMux I__4564 (
            .O(N__19866),
            .I(N__19857));
    LocalMux I__4563 (
            .O(N__19863),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__4562 (
            .O(N__19860),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__4561 (
            .O(N__19857),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__4560 (
            .O(N__19850),
            .I(N__19847));
    LocalMux I__4559 (
            .O(N__19847),
            .I(N__19844));
    Span4Mux_h I__4558 (
            .O(N__19844),
            .I(N__19840));
    InMux I__4557 (
            .O(N__19843),
            .I(N__19837));
    Span4Mux_v I__4556 (
            .O(N__19840),
            .I(N__19834));
    LocalMux I__4555 (
            .O(N__19837),
            .I(N__19831));
    Odrv4 I__4554 (
            .O(N__19834),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    Odrv12 I__4553 (
            .O(N__19831),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__4552 (
            .O(N__19826),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__4551 (
            .O(N__19823),
            .I(N__19818));
    InMux I__4550 (
            .O(N__19822),
            .I(N__19815));
    InMux I__4549 (
            .O(N__19821),
            .I(N__19812));
    InMux I__4548 (
            .O(N__19818),
            .I(N__19809));
    LocalMux I__4547 (
            .O(N__19815),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__4546 (
            .O(N__19812),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__4545 (
            .O(N__19809),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__4544 (
            .O(N__19802),
            .I(N__19798));
    CascadeMux I__4543 (
            .O(N__19801),
            .I(N__19794));
    LocalMux I__4542 (
            .O(N__19798),
            .I(N__19791));
    InMux I__4541 (
            .O(N__19797),
            .I(N__19788));
    InMux I__4540 (
            .O(N__19794),
            .I(N__19785));
    Span4Mux_v I__4539 (
            .O(N__19791),
            .I(N__19778));
    LocalMux I__4538 (
            .O(N__19788),
            .I(N__19778));
    LocalMux I__4537 (
            .O(N__19785),
            .I(N__19778));
    Span4Mux_h I__4536 (
            .O(N__19778),
            .I(N__19775));
    Odrv4 I__4535 (
            .O(N__19775),
            .I(\delay_measurement_inst.elapsed_time_tr_9 ));
    InMux I__4534 (
            .O(N__19772),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__4533 (
            .O(N__19769),
            .I(N__19764));
    InMux I__4532 (
            .O(N__19768),
            .I(N__19761));
    InMux I__4531 (
            .O(N__19767),
            .I(N__19758));
    InMux I__4530 (
            .O(N__19764),
            .I(N__19755));
    LocalMux I__4529 (
            .O(N__19761),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__4528 (
            .O(N__19758),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__4527 (
            .O(N__19755),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__4526 (
            .O(N__19748),
            .I(N__19745));
    LocalMux I__4525 (
            .O(N__19745),
            .I(N__19741));
    InMux I__4524 (
            .O(N__19744),
            .I(N__19738));
    Span4Mux_v I__4523 (
            .O(N__19741),
            .I(N__19733));
    LocalMux I__4522 (
            .O(N__19738),
            .I(N__19733));
    Span4Mux_h I__4521 (
            .O(N__19733),
            .I(N__19730));
    Odrv4 I__4520 (
            .O(N__19730),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__4519 (
            .O(N__19727),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__4518 (
            .O(N__19724),
            .I(N__19719));
    InMux I__4517 (
            .O(N__19723),
            .I(N__19716));
    InMux I__4516 (
            .O(N__19722),
            .I(N__19713));
    InMux I__4515 (
            .O(N__19719),
            .I(N__19710));
    LocalMux I__4514 (
            .O(N__19716),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__4513 (
            .O(N__19713),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__4512 (
            .O(N__19710),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__4511 (
            .O(N__19703),
            .I(N__19699));
    InMux I__4510 (
            .O(N__19702),
            .I(N__19696));
    LocalMux I__4509 (
            .O(N__19699),
            .I(N__19693));
    LocalMux I__4508 (
            .O(N__19696),
            .I(N__19690));
    Span4Mux_h I__4507 (
            .O(N__19693),
            .I(N__19687));
    Odrv12 I__4506 (
            .O(N__19690),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    Odrv4 I__4505 (
            .O(N__19687),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__4504 (
            .O(N__19682),
            .I(bfn_13_20_0_));
    CascadeMux I__4503 (
            .O(N__19679),
            .I(N__19674));
    InMux I__4502 (
            .O(N__19678),
            .I(N__19671));
    InMux I__4501 (
            .O(N__19677),
            .I(N__19668));
    InMux I__4500 (
            .O(N__19674),
            .I(N__19665));
    LocalMux I__4499 (
            .O(N__19671),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__4498 (
            .O(N__19668),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__4497 (
            .O(N__19665),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__4496 (
            .O(N__19658),
            .I(N__19654));
    InMux I__4495 (
            .O(N__19657),
            .I(N__19651));
    LocalMux I__4494 (
            .O(N__19654),
            .I(N__19648));
    LocalMux I__4493 (
            .O(N__19651),
            .I(N__19645));
    Span4Mux_h I__4492 (
            .O(N__19648),
            .I(N__19642));
    Odrv12 I__4491 (
            .O(N__19645),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    Odrv4 I__4490 (
            .O(N__19642),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__4489 (
            .O(N__19637),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__4488 (
            .O(N__19634),
            .I(N__19629));
    InMux I__4487 (
            .O(N__19633),
            .I(N__19626));
    InMux I__4486 (
            .O(N__19632),
            .I(N__19623));
    InMux I__4485 (
            .O(N__19629),
            .I(N__19620));
    LocalMux I__4484 (
            .O(N__19626),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__4483 (
            .O(N__19623),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__4482 (
            .O(N__19620),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    CascadeMux I__4481 (
            .O(N__19613),
            .I(N__19609));
    InMux I__4480 (
            .O(N__19612),
            .I(N__19606));
    InMux I__4479 (
            .O(N__19609),
            .I(N__19603));
    LocalMux I__4478 (
            .O(N__19606),
            .I(N__19600));
    LocalMux I__4477 (
            .O(N__19603),
            .I(N__19597));
    Span4Mux_h I__4476 (
            .O(N__19600),
            .I(N__19594));
    Span4Mux_h I__4475 (
            .O(N__19597),
            .I(N__19591));
    Odrv4 I__4474 (
            .O(N__19594),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    Odrv4 I__4473 (
            .O(N__19591),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    InMux I__4472 (
            .O(N__19586),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__4471 (
            .O(N__19583),
            .I(N__19578));
    InMux I__4470 (
            .O(N__19582),
            .I(N__19575));
    InMux I__4469 (
            .O(N__19581),
            .I(N__19572));
    InMux I__4468 (
            .O(N__19578),
            .I(N__19569));
    LocalMux I__4467 (
            .O(N__19575),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__4466 (
            .O(N__19572),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__4465 (
            .O(N__19569),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    CascadeMux I__4464 (
            .O(N__19562),
            .I(N__19559));
    InMux I__4463 (
            .O(N__19559),
            .I(N__19553));
    InMux I__4462 (
            .O(N__19558),
            .I(N__19548));
    InMux I__4461 (
            .O(N__19557),
            .I(N__19548));
    InMux I__4460 (
            .O(N__19556),
            .I(N__19545));
    LocalMux I__4459 (
            .O(N__19553),
            .I(N__19540));
    LocalMux I__4458 (
            .O(N__19548),
            .I(N__19540));
    LocalMux I__4457 (
            .O(N__19545),
            .I(N__19537));
    Span4Mux_h I__4456 (
            .O(N__19540),
            .I(N__19534));
    Odrv12 I__4455 (
            .O(N__19537),
            .I(\delay_measurement_inst.elapsed_time_tr_14 ));
    Odrv4 I__4454 (
            .O(N__19534),
            .I(\delay_measurement_inst.elapsed_time_tr_14 ));
    InMux I__4453 (
            .O(N__19529),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__4452 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__4451 (
            .O(N__19523),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    InMux I__4450 (
            .O(N__19520),
            .I(N__19516));
    InMux I__4449 (
            .O(N__19519),
            .I(N__19513));
    LocalMux I__4448 (
            .O(N__19516),
            .I(N__19510));
    LocalMux I__4447 (
            .O(N__19513),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__4446 (
            .O(N__19510),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__4445 (
            .O(N__19505),
            .I(N__19501));
    CascadeMux I__4444 (
            .O(N__19504),
            .I(N__19497));
    LocalMux I__4443 (
            .O(N__19501),
            .I(N__19494));
    InMux I__4442 (
            .O(N__19500),
            .I(N__19491));
    InMux I__4441 (
            .O(N__19497),
            .I(N__19488));
    Span4Mux_v I__4440 (
            .O(N__19494),
            .I(N__19485));
    LocalMux I__4439 (
            .O(N__19491),
            .I(N__19481));
    LocalMux I__4438 (
            .O(N__19488),
            .I(N__19476));
    Span4Mux_h I__4437 (
            .O(N__19485),
            .I(N__19476));
    InMux I__4436 (
            .O(N__19484),
            .I(N__19473));
    Span4Mux_v I__4435 (
            .O(N__19481),
            .I(N__19470));
    Odrv4 I__4434 (
            .O(N__19476),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__4433 (
            .O(N__19473),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__4432 (
            .O(N__19470),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    CascadeMux I__4431 (
            .O(N__19463),
            .I(N__19452));
    CascadeMux I__4430 (
            .O(N__19462),
            .I(N__19449));
    CascadeMux I__4429 (
            .O(N__19461),
            .I(N__19446));
    CascadeMux I__4428 (
            .O(N__19460),
            .I(N__19442));
    InMux I__4427 (
            .O(N__19459),
            .I(N__19439));
    InMux I__4426 (
            .O(N__19458),
            .I(N__19417));
    InMux I__4425 (
            .O(N__19457),
            .I(N__19417));
    InMux I__4424 (
            .O(N__19456),
            .I(N__19417));
    InMux I__4423 (
            .O(N__19455),
            .I(N__19417));
    InMux I__4422 (
            .O(N__19452),
            .I(N__19417));
    InMux I__4421 (
            .O(N__19449),
            .I(N__19417));
    InMux I__4420 (
            .O(N__19446),
            .I(N__19417));
    InMux I__4419 (
            .O(N__19445),
            .I(N__19414));
    InMux I__4418 (
            .O(N__19442),
            .I(N__19411));
    LocalMux I__4417 (
            .O(N__19439),
            .I(N__19408));
    CascadeMux I__4416 (
            .O(N__19438),
            .I(N__19404));
    CascadeMux I__4415 (
            .O(N__19437),
            .I(N__19401));
    CascadeMux I__4414 (
            .O(N__19436),
            .I(N__19398));
    CascadeMux I__4413 (
            .O(N__19435),
            .I(N__19395));
    CascadeMux I__4412 (
            .O(N__19434),
            .I(N__19389));
    CascadeMux I__4411 (
            .O(N__19433),
            .I(N__19386));
    CascadeMux I__4410 (
            .O(N__19432),
            .I(N__19383));
    LocalMux I__4409 (
            .O(N__19417),
            .I(N__19378));
    LocalMux I__4408 (
            .O(N__19414),
            .I(N__19375));
    LocalMux I__4407 (
            .O(N__19411),
            .I(N__19370));
    Span4Mux_v I__4406 (
            .O(N__19408),
            .I(N__19370));
    InMux I__4405 (
            .O(N__19407),
            .I(N__19353));
    InMux I__4404 (
            .O(N__19404),
            .I(N__19353));
    InMux I__4403 (
            .O(N__19401),
            .I(N__19353));
    InMux I__4402 (
            .O(N__19398),
            .I(N__19353));
    InMux I__4401 (
            .O(N__19395),
            .I(N__19353));
    InMux I__4400 (
            .O(N__19394),
            .I(N__19353));
    InMux I__4399 (
            .O(N__19393),
            .I(N__19353));
    InMux I__4398 (
            .O(N__19392),
            .I(N__19353));
    InMux I__4397 (
            .O(N__19389),
            .I(N__19342));
    InMux I__4396 (
            .O(N__19386),
            .I(N__19342));
    InMux I__4395 (
            .O(N__19383),
            .I(N__19342));
    InMux I__4394 (
            .O(N__19382),
            .I(N__19342));
    InMux I__4393 (
            .O(N__19381),
            .I(N__19342));
    Span4Mux_h I__4392 (
            .O(N__19378),
            .I(N__19339));
    Span4Mux_v I__4391 (
            .O(N__19375),
            .I(N__19334));
    Span4Mux_h I__4390 (
            .O(N__19370),
            .I(N__19334));
    LocalMux I__4389 (
            .O(N__19353),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__4388 (
            .O(N__19342),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__4387 (
            .O(N__19339),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__4386 (
            .O(N__19334),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    InMux I__4385 (
            .O(N__19325),
            .I(N__19322));
    LocalMux I__4384 (
            .O(N__19322),
            .I(N__19319));
    Span4Mux_v I__4383 (
            .O(N__19319),
            .I(N__19316));
    Odrv4 I__4382 (
            .O(N__19316),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__4381 (
            .O(N__19313),
            .I(N__19310));
    LocalMux I__4380 (
            .O(N__19310),
            .I(\phase_controller_inst1.N_112 ));
    InMux I__4379 (
            .O(N__19307),
            .I(N__19286));
    InMux I__4378 (
            .O(N__19306),
            .I(N__19286));
    InMux I__4377 (
            .O(N__19305),
            .I(N__19286));
    InMux I__4376 (
            .O(N__19304),
            .I(N__19286));
    InMux I__4375 (
            .O(N__19303),
            .I(N__19286));
    InMux I__4374 (
            .O(N__19302),
            .I(N__19286));
    InMux I__4373 (
            .O(N__19301),
            .I(N__19286));
    LocalMux I__4372 (
            .O(N__19286),
            .I(N__19269));
    InMux I__4371 (
            .O(N__19285),
            .I(N__19260));
    InMux I__4370 (
            .O(N__19284),
            .I(N__19260));
    InMux I__4369 (
            .O(N__19283),
            .I(N__19260));
    InMux I__4368 (
            .O(N__19282),
            .I(N__19260));
    InMux I__4367 (
            .O(N__19281),
            .I(N__19257));
    InMux I__4366 (
            .O(N__19280),
            .I(N__19240));
    InMux I__4365 (
            .O(N__19279),
            .I(N__19240));
    InMux I__4364 (
            .O(N__19278),
            .I(N__19240));
    InMux I__4363 (
            .O(N__19277),
            .I(N__19240));
    InMux I__4362 (
            .O(N__19276),
            .I(N__19240));
    InMux I__4361 (
            .O(N__19275),
            .I(N__19240));
    InMux I__4360 (
            .O(N__19274),
            .I(N__19240));
    InMux I__4359 (
            .O(N__19273),
            .I(N__19240));
    CascadeMux I__4358 (
            .O(N__19272),
            .I(N__19235));
    Span4Mux_h I__4357 (
            .O(N__19269),
            .I(N__19232));
    LocalMux I__4356 (
            .O(N__19260),
            .I(N__19227));
    LocalMux I__4355 (
            .O(N__19257),
            .I(N__19227));
    LocalMux I__4354 (
            .O(N__19240),
            .I(N__19224));
    InMux I__4353 (
            .O(N__19239),
            .I(N__19220));
    InMux I__4352 (
            .O(N__19238),
            .I(N__19217));
    InMux I__4351 (
            .O(N__19235),
            .I(N__19214));
    Span4Mux_v I__4350 (
            .O(N__19232),
            .I(N__19211));
    Span4Mux_h I__4349 (
            .O(N__19227),
            .I(N__19208));
    Span4Mux_h I__4348 (
            .O(N__19224),
            .I(N__19205));
    InMux I__4347 (
            .O(N__19223),
            .I(N__19202));
    LocalMux I__4346 (
            .O(N__19220),
            .I(N__19197));
    LocalMux I__4345 (
            .O(N__19217),
            .I(N__19197));
    LocalMux I__4344 (
            .O(N__19214),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__4343 (
            .O(N__19211),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__4342 (
            .O(N__19208),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__4341 (
            .O(N__19205),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__4340 (
            .O(N__19202),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__4339 (
            .O(N__19197),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__4338 (
            .O(N__19184),
            .I(N__19179));
    InMux I__4337 (
            .O(N__19183),
            .I(N__19176));
    InMux I__4336 (
            .O(N__19182),
            .I(N__19173));
    LocalMux I__4335 (
            .O(N__19179),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__4334 (
            .O(N__19176),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__4333 (
            .O(N__19173),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__4332 (
            .O(N__19166),
            .I(N__19162));
    InMux I__4331 (
            .O(N__19165),
            .I(N__19159));
    LocalMux I__4330 (
            .O(N__19162),
            .I(N__19156));
    LocalMux I__4329 (
            .O(N__19159),
            .I(N__19153));
    Span4Mux_h I__4328 (
            .O(N__19156),
            .I(N__19150));
    Span4Mux_h I__4327 (
            .O(N__19153),
            .I(N__19147));
    Odrv4 I__4326 (
            .O(N__19150),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    Odrv4 I__4325 (
            .O(N__19147),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    InMux I__4324 (
            .O(N__19142),
            .I(N__19137));
    InMux I__4323 (
            .O(N__19141),
            .I(N__19134));
    InMux I__4322 (
            .O(N__19140),
            .I(N__19131));
    LocalMux I__4321 (
            .O(N__19137),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__4320 (
            .O(N__19134),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__4319 (
            .O(N__19131),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    CascadeMux I__4318 (
            .O(N__19124),
            .I(N__19121));
    InMux I__4317 (
            .O(N__19121),
            .I(N__19117));
    InMux I__4316 (
            .O(N__19120),
            .I(N__19114));
    LocalMux I__4315 (
            .O(N__19117),
            .I(N__19111));
    LocalMux I__4314 (
            .O(N__19114),
            .I(N__19108));
    Span4Mux_h I__4313 (
            .O(N__19111),
            .I(N__19105));
    Span4Mux_h I__4312 (
            .O(N__19108),
            .I(N__19102));
    Odrv4 I__4311 (
            .O(N__19105),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    Odrv4 I__4310 (
            .O(N__19102),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    InMux I__4309 (
            .O(N__19097),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__4308 (
            .O(N__19094),
            .I(N__19089));
    InMux I__4307 (
            .O(N__19093),
            .I(N__19086));
    InMux I__4306 (
            .O(N__19092),
            .I(N__19083));
    InMux I__4305 (
            .O(N__19089),
            .I(N__19080));
    LocalMux I__4304 (
            .O(N__19086),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__4303 (
            .O(N__19083),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__4302 (
            .O(N__19080),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__4301 (
            .O(N__19073),
            .I(N__19069));
    InMux I__4300 (
            .O(N__19072),
            .I(N__19066));
    LocalMux I__4299 (
            .O(N__19069),
            .I(N__19063));
    LocalMux I__4298 (
            .O(N__19066),
            .I(N__19060));
    Span4Mux_h I__4297 (
            .O(N__19063),
            .I(N__19057));
    Span4Mux_v I__4296 (
            .O(N__19060),
            .I(N__19054));
    Odrv4 I__4295 (
            .O(N__19057),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    Odrv4 I__4294 (
            .O(N__19054),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__4293 (
            .O(N__19049),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__4292 (
            .O(N__19046),
            .I(N__19041));
    InMux I__4291 (
            .O(N__19045),
            .I(N__19038));
    InMux I__4290 (
            .O(N__19044),
            .I(N__19035));
    InMux I__4289 (
            .O(N__19041),
            .I(N__19032));
    LocalMux I__4288 (
            .O(N__19038),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__4287 (
            .O(N__19035),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__4286 (
            .O(N__19032),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__4285 (
            .O(N__19025),
            .I(N__19022));
    LocalMux I__4284 (
            .O(N__19022),
            .I(N__19018));
    InMux I__4283 (
            .O(N__19021),
            .I(N__19015));
    Span4Mux_h I__4282 (
            .O(N__19018),
            .I(N__19012));
    LocalMux I__4281 (
            .O(N__19015),
            .I(N__19009));
    Odrv4 I__4280 (
            .O(N__19012),
            .I(\delay_measurement_inst.elapsed_time_tr_6 ));
    Odrv12 I__4279 (
            .O(N__19009),
            .I(\delay_measurement_inst.elapsed_time_tr_6 ));
    InMux I__4278 (
            .O(N__19004),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__4277 (
            .O(N__19001),
            .I(N__18996));
    InMux I__4276 (
            .O(N__19000),
            .I(N__18993));
    InMux I__4275 (
            .O(N__18999),
            .I(N__18990));
    InMux I__4274 (
            .O(N__18996),
            .I(N__18987));
    LocalMux I__4273 (
            .O(N__18993),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__4272 (
            .O(N__18990),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__4271 (
            .O(N__18987),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__4270 (
            .O(N__18980),
            .I(N__18977));
    LocalMux I__4269 (
            .O(N__18977),
            .I(N__18973));
    InMux I__4268 (
            .O(N__18976),
            .I(N__18970));
    Span4Mux_h I__4267 (
            .O(N__18973),
            .I(N__18963));
    LocalMux I__4266 (
            .O(N__18970),
            .I(N__18963));
    InMux I__4265 (
            .O(N__18969),
            .I(N__18960));
    InMux I__4264 (
            .O(N__18968),
            .I(N__18957));
    Odrv4 I__4263 (
            .O(N__18963),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__4262 (
            .O(N__18960),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__4261 (
            .O(N__18957),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__4260 (
            .O(N__18950),
            .I(N__18947));
    LocalMux I__4259 (
            .O(N__18947),
            .I(N__18944));
    Span4Mux_s2_v I__4258 (
            .O(N__18944),
            .I(N__18941));
    Odrv4 I__4257 (
            .O(N__18941),
            .I(s2_phy_c));
    InMux I__4256 (
            .O(N__18938),
            .I(N__18933));
    CascadeMux I__4255 (
            .O(N__18937),
            .I(N__18930));
    CascadeMux I__4254 (
            .O(N__18936),
            .I(N__18927));
    LocalMux I__4253 (
            .O(N__18933),
            .I(N__18924));
    InMux I__4252 (
            .O(N__18930),
            .I(N__18921));
    InMux I__4251 (
            .O(N__18927),
            .I(N__18917));
    Span4Mux_v I__4250 (
            .O(N__18924),
            .I(N__18912));
    LocalMux I__4249 (
            .O(N__18921),
            .I(N__18912));
    InMux I__4248 (
            .O(N__18920),
            .I(N__18909));
    LocalMux I__4247 (
            .O(N__18917),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    Odrv4 I__4246 (
            .O(N__18912),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__4245 (
            .O(N__18909),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    IoInMux I__4244 (
            .O(N__18902),
            .I(N__18899));
    LocalMux I__4243 (
            .O(N__18899),
            .I(N__18896));
    Span4Mux_s1_v I__4242 (
            .O(N__18896),
            .I(N__18893));
    Odrv4 I__4241 (
            .O(N__18893),
            .I(s1_phy_c));
    IoInMux I__4240 (
            .O(N__18890),
            .I(N__18887));
    LocalMux I__4239 (
            .O(N__18887),
            .I(N__18884));
    Span4Mux_s0_v I__4238 (
            .O(N__18884),
            .I(N__18881));
    Odrv4 I__4237 (
            .O(N__18881),
            .I(\pll_inst.red_c_i ));
    InMux I__4236 (
            .O(N__18878),
            .I(N__18875));
    LocalMux I__4235 (
            .O(N__18875),
            .I(N__18872));
    Span4Mux_h I__4234 (
            .O(N__18872),
            .I(N__18869));
    Span4Mux_v I__4233 (
            .O(N__18869),
            .I(N__18866));
    Odrv4 I__4232 (
            .O(N__18866),
            .I(delay_hc_input_c));
    InMux I__4231 (
            .O(N__18863),
            .I(N__18860));
    LocalMux I__4230 (
            .O(N__18860),
            .I(delay_hc_d1));
    InMux I__4229 (
            .O(N__18857),
            .I(N__18854));
    LocalMux I__4228 (
            .O(N__18854),
            .I(N__18851));
    Odrv12 I__4227 (
            .O(N__18851),
            .I(\delay_measurement_inst.tr_syncZ0Z_0 ));
    InMux I__4226 (
            .O(N__18848),
            .I(N__18844));
    InMux I__4225 (
            .O(N__18847),
            .I(N__18841));
    LocalMux I__4224 (
            .O(N__18844),
            .I(N__18836));
    LocalMux I__4223 (
            .O(N__18841),
            .I(N__18836));
    Span4Mux_h I__4222 (
            .O(N__18836),
            .I(N__18833));
    Odrv4 I__4221 (
            .O(N__18833),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__4220 (
            .O(N__18830),
            .I(N__18826));
    InMux I__4219 (
            .O(N__18829),
            .I(N__18823));
    LocalMux I__4218 (
            .O(N__18826),
            .I(N__18817));
    LocalMux I__4217 (
            .O(N__18823),
            .I(N__18817));
    InMux I__4216 (
            .O(N__18822),
            .I(N__18814));
    Span4Mux_v I__4215 (
            .O(N__18817),
            .I(N__18811));
    LocalMux I__4214 (
            .O(N__18814),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__4213 (
            .O(N__18811),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__4212 (
            .O(N__18806),
            .I(N__18800));
    InMux I__4211 (
            .O(N__18805),
            .I(N__18795));
    InMux I__4210 (
            .O(N__18804),
            .I(N__18795));
    InMux I__4209 (
            .O(N__18803),
            .I(N__18792));
    LocalMux I__4208 (
            .O(N__18800),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__4207 (
            .O(N__18795),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__4206 (
            .O(N__18792),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    IoInMux I__4205 (
            .O(N__18785),
            .I(N__18782));
    LocalMux I__4204 (
            .O(N__18782),
            .I(N__18779));
    Span12Mux_s8_v I__4203 (
            .O(N__18779),
            .I(N__18776));
    Odrv12 I__4202 (
            .O(N__18776),
            .I(\delay_measurement_inst.delay_hc_timer.N_178_i ));
    CEMux I__4201 (
            .O(N__18773),
            .I(N__18769));
    CEMux I__4200 (
            .O(N__18772),
            .I(N__18766));
    LocalMux I__4199 (
            .O(N__18769),
            .I(N__18762));
    LocalMux I__4198 (
            .O(N__18766),
            .I(N__18759));
    CEMux I__4197 (
            .O(N__18765),
            .I(N__18756));
    Span4Mux_h I__4196 (
            .O(N__18762),
            .I(N__18753));
    Span4Mux_h I__4195 (
            .O(N__18759),
            .I(N__18750));
    LocalMux I__4194 (
            .O(N__18756),
            .I(N__18747));
    Odrv4 I__4193 (
            .O(N__18753),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1 ));
    Odrv4 I__4192 (
            .O(N__18750),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1 ));
    Odrv12 I__4191 (
            .O(N__18747),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1 ));
    InMux I__4190 (
            .O(N__18740),
            .I(bfn_12_21_0_));
    InMux I__4189 (
            .O(N__18737),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__4188 (
            .O(N__18734),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__4187 (
            .O(N__18731),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__4186 (
            .O(N__18728),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__4185 (
            .O(N__18725),
            .I(N__18687));
    InMux I__4184 (
            .O(N__18724),
            .I(N__18687));
    InMux I__4183 (
            .O(N__18723),
            .I(N__18687));
    InMux I__4182 (
            .O(N__18722),
            .I(N__18687));
    InMux I__4181 (
            .O(N__18721),
            .I(N__18678));
    InMux I__4180 (
            .O(N__18720),
            .I(N__18678));
    InMux I__4179 (
            .O(N__18719),
            .I(N__18678));
    InMux I__4178 (
            .O(N__18718),
            .I(N__18678));
    InMux I__4177 (
            .O(N__18717),
            .I(N__18669));
    InMux I__4176 (
            .O(N__18716),
            .I(N__18669));
    InMux I__4175 (
            .O(N__18715),
            .I(N__18669));
    InMux I__4174 (
            .O(N__18714),
            .I(N__18669));
    InMux I__4173 (
            .O(N__18713),
            .I(N__18664));
    InMux I__4172 (
            .O(N__18712),
            .I(N__18664));
    InMux I__4171 (
            .O(N__18711),
            .I(N__18655));
    InMux I__4170 (
            .O(N__18710),
            .I(N__18655));
    InMux I__4169 (
            .O(N__18709),
            .I(N__18655));
    InMux I__4168 (
            .O(N__18708),
            .I(N__18655));
    InMux I__4167 (
            .O(N__18707),
            .I(N__18646));
    InMux I__4166 (
            .O(N__18706),
            .I(N__18646));
    InMux I__4165 (
            .O(N__18705),
            .I(N__18646));
    InMux I__4164 (
            .O(N__18704),
            .I(N__18646));
    InMux I__4163 (
            .O(N__18703),
            .I(N__18637));
    InMux I__4162 (
            .O(N__18702),
            .I(N__18637));
    InMux I__4161 (
            .O(N__18701),
            .I(N__18637));
    InMux I__4160 (
            .O(N__18700),
            .I(N__18637));
    InMux I__4159 (
            .O(N__18699),
            .I(N__18628));
    InMux I__4158 (
            .O(N__18698),
            .I(N__18628));
    InMux I__4157 (
            .O(N__18697),
            .I(N__18628));
    InMux I__4156 (
            .O(N__18696),
            .I(N__18628));
    LocalMux I__4155 (
            .O(N__18687),
            .I(N__18621));
    LocalMux I__4154 (
            .O(N__18678),
            .I(N__18621));
    LocalMux I__4153 (
            .O(N__18669),
            .I(N__18621));
    LocalMux I__4152 (
            .O(N__18664),
            .I(N__18610));
    LocalMux I__4151 (
            .O(N__18655),
            .I(N__18610));
    LocalMux I__4150 (
            .O(N__18646),
            .I(N__18610));
    LocalMux I__4149 (
            .O(N__18637),
            .I(N__18610));
    LocalMux I__4148 (
            .O(N__18628),
            .I(N__18610));
    Span4Mux_v I__4147 (
            .O(N__18621),
            .I(N__18605));
    Span4Mux_v I__4146 (
            .O(N__18610),
            .I(N__18605));
    Span4Mux_v I__4145 (
            .O(N__18605),
            .I(N__18602));
    Odrv4 I__4144 (
            .O(N__18602),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__4143 (
            .O(N__18599),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__4142 (
            .O(N__18596),
            .I(N__18584));
    CEMux I__4141 (
            .O(N__18595),
            .I(N__18584));
    CEMux I__4140 (
            .O(N__18594),
            .I(N__18584));
    CEMux I__4139 (
            .O(N__18593),
            .I(N__18584));
    GlobalMux I__4138 (
            .O(N__18584),
            .I(N__18581));
    gio2CtrlBuf I__4137 (
            .O(N__18581),
            .I(\delay_measurement_inst.delay_tr_timer.N_181_i_g ));
    InMux I__4136 (
            .O(N__18578),
            .I(N__18573));
    InMux I__4135 (
            .O(N__18577),
            .I(N__18570));
    InMux I__4134 (
            .O(N__18576),
            .I(N__18567));
    LocalMux I__4133 (
            .O(N__18573),
            .I(N__18560));
    LocalMux I__4132 (
            .O(N__18570),
            .I(N__18560));
    LocalMux I__4131 (
            .O(N__18567),
            .I(N__18560));
    Span12Mux_s11_v I__4130 (
            .O(N__18560),
            .I(N__18557));
    Odrv12 I__4129 (
            .O(N__18557),
            .I(il_max_comp1_D2));
    InMux I__4128 (
            .O(N__18554),
            .I(N__18551));
    LocalMux I__4127 (
            .O(N__18551),
            .I(N__18548));
    Span4Mux_h I__4126 (
            .O(N__18548),
            .I(N__18544));
    InMux I__4125 (
            .O(N__18547),
            .I(N__18541));
    Odrv4 I__4124 (
            .O(N__18544),
            .I(\phase_controller_inst1.N_108 ));
    LocalMux I__4123 (
            .O(N__18541),
            .I(\phase_controller_inst1.N_108 ));
    InMux I__4122 (
            .O(N__18536),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__4121 (
            .O(N__18533),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__4120 (
            .O(N__18530),
            .I(bfn_12_20_0_));
    InMux I__4119 (
            .O(N__18527),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__4118 (
            .O(N__18524),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__4117 (
            .O(N__18521),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__4116 (
            .O(N__18518),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__4115 (
            .O(N__18515),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__4114 (
            .O(N__18512),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__4113 (
            .O(N__18509),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__4112 (
            .O(N__18506),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__4111 (
            .O(N__18503),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__4110 (
            .O(N__18500),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__4109 (
            .O(N__18497),
            .I(bfn_12_19_0_));
    InMux I__4108 (
            .O(N__18494),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__4107 (
            .O(N__18491),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__4106 (
            .O(N__18488),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__4105 (
            .O(N__18485),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__4104 (
            .O(N__18482),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__4103 (
            .O(N__18479),
            .I(N__18475));
    InMux I__4102 (
            .O(N__18478),
            .I(N__18472));
    LocalMux I__4101 (
            .O(N__18475),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__4100 (
            .O(N__18472),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__4099 (
            .O(N__18467),
            .I(N__18464));
    LocalMux I__4098 (
            .O(N__18464),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__4097 (
            .O(N__18461),
            .I(bfn_12_17_0_));
    InMux I__4096 (
            .O(N__18458),
            .I(N__18454));
    InMux I__4095 (
            .O(N__18457),
            .I(N__18451));
    LocalMux I__4094 (
            .O(N__18454),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__4093 (
            .O(N__18451),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__4092 (
            .O(N__18446),
            .I(N__18443));
    LocalMux I__4091 (
            .O(N__18443),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    InMux I__4090 (
            .O(N__18440),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__4089 (
            .O(N__18437),
            .I(N__18433));
    InMux I__4088 (
            .O(N__18436),
            .I(N__18430));
    LocalMux I__4087 (
            .O(N__18433),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__4086 (
            .O(N__18430),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__4085 (
            .O(N__18425),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__4084 (
            .O(N__18422),
            .I(N__18419));
    LocalMux I__4083 (
            .O(N__18419),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    InMux I__4082 (
            .O(N__18416),
            .I(bfn_12_18_0_));
    InMux I__4081 (
            .O(N__18413),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__4080 (
            .O(N__18410),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__4079 (
            .O(N__18407),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__4078 (
            .O(N__18404),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__4077 (
            .O(N__18401),
            .I(N__18397));
    InMux I__4076 (
            .O(N__18400),
            .I(N__18394));
    LocalMux I__4075 (
            .O(N__18397),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__4074 (
            .O(N__18394),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__4073 (
            .O(N__18389),
            .I(N__18386));
    InMux I__4072 (
            .O(N__18386),
            .I(N__18383));
    LocalMux I__4071 (
            .O(N__18383),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__4070 (
            .O(N__18380),
            .I(bfn_12_16_0_));
    InMux I__4069 (
            .O(N__18377),
            .I(N__18373));
    InMux I__4068 (
            .O(N__18376),
            .I(N__18370));
    LocalMux I__4067 (
            .O(N__18373),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__4066 (
            .O(N__18370),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__4065 (
            .O(N__18365),
            .I(N__18362));
    LocalMux I__4064 (
            .O(N__18362),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__4063 (
            .O(N__18359),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__4062 (
            .O(N__18356),
            .I(N__18352));
    InMux I__4061 (
            .O(N__18355),
            .I(N__18349));
    LocalMux I__4060 (
            .O(N__18352),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__4059 (
            .O(N__18349),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__4058 (
            .O(N__18344),
            .I(N__18341));
    LocalMux I__4057 (
            .O(N__18341),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    InMux I__4056 (
            .O(N__18338),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__4055 (
            .O(N__18335),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__4054 (
            .O(N__18332),
            .I(N__18328));
    InMux I__4053 (
            .O(N__18331),
            .I(N__18325));
    LocalMux I__4052 (
            .O(N__18328),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__4051 (
            .O(N__18325),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__4050 (
            .O(N__18320),
            .I(N__18317));
    LocalMux I__4049 (
            .O(N__18317),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__4048 (
            .O(N__18314),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__4047 (
            .O(N__18311),
            .I(N__18307));
    InMux I__4046 (
            .O(N__18310),
            .I(N__18304));
    LocalMux I__4045 (
            .O(N__18307),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__4044 (
            .O(N__18304),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__4043 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__4042 (
            .O(N__18296),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__4041 (
            .O(N__18293),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__4040 (
            .O(N__18290),
            .I(N__18286));
    InMux I__4039 (
            .O(N__18289),
            .I(N__18283));
    LocalMux I__4038 (
            .O(N__18286),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__4037 (
            .O(N__18283),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__4036 (
            .O(N__18278),
            .I(N__18275));
    LocalMux I__4035 (
            .O(N__18275),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    InMux I__4034 (
            .O(N__18272),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__4033 (
            .O(N__18269),
            .I(N__18265));
    InMux I__4032 (
            .O(N__18268),
            .I(N__18262));
    LocalMux I__4031 (
            .O(N__18265),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__4030 (
            .O(N__18262),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__4029 (
            .O(N__18257),
            .I(N__18254));
    LocalMux I__4028 (
            .O(N__18254),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    InMux I__4027 (
            .O(N__18251),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__4026 (
            .O(N__18248),
            .I(N__18243));
    InMux I__4025 (
            .O(N__18247),
            .I(N__18240));
    InMux I__4024 (
            .O(N__18246),
            .I(N__18237));
    LocalMux I__4023 (
            .O(N__18243),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__4022 (
            .O(N__18240),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__4021 (
            .O(N__18237),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__4020 (
            .O(N__18230),
            .I(N__18227));
    InMux I__4019 (
            .O(N__18227),
            .I(N__18224));
    LocalMux I__4018 (
            .O(N__18224),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    InMux I__4017 (
            .O(N__18221),
            .I(N__18217));
    InMux I__4016 (
            .O(N__18220),
            .I(N__18214));
    LocalMux I__4015 (
            .O(N__18217),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__4014 (
            .O(N__18214),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__4013 (
            .O(N__18209),
            .I(N__18206));
    InMux I__4012 (
            .O(N__18206),
            .I(N__18203));
    LocalMux I__4011 (
            .O(N__18203),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__4010 (
            .O(N__18200),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__4009 (
            .O(N__18197),
            .I(N__18193));
    InMux I__4008 (
            .O(N__18196),
            .I(N__18190));
    LocalMux I__4007 (
            .O(N__18193),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__4006 (
            .O(N__18190),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__4005 (
            .O(N__18185),
            .I(N__18182));
    InMux I__4004 (
            .O(N__18182),
            .I(N__18179));
    LocalMux I__4003 (
            .O(N__18179),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0 ));
    CascadeMux I__4002 (
            .O(N__18176),
            .I(N__18173));
    InMux I__4001 (
            .O(N__18173),
            .I(N__18170));
    LocalMux I__4000 (
            .O(N__18170),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    InMux I__3999 (
            .O(N__18167),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__3998 (
            .O(N__18164),
            .I(N__18160));
    InMux I__3997 (
            .O(N__18163),
            .I(N__18157));
    LocalMux I__3996 (
            .O(N__18160),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__3995 (
            .O(N__18157),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__3994 (
            .O(N__18152),
            .I(N__18149));
    LocalMux I__3993 (
            .O(N__18149),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__3992 (
            .O(N__18146),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    CascadeMux I__3991 (
            .O(N__18143),
            .I(N__18140));
    InMux I__3990 (
            .O(N__18140),
            .I(N__18136));
    InMux I__3989 (
            .O(N__18139),
            .I(N__18133));
    LocalMux I__3988 (
            .O(N__18136),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__3987 (
            .O(N__18133),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__3986 (
            .O(N__18128),
            .I(N__18125));
    InMux I__3985 (
            .O(N__18125),
            .I(N__18122));
    LocalMux I__3984 (
            .O(N__18122),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__3983 (
            .O(N__18119),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    CascadeMux I__3982 (
            .O(N__18116),
            .I(N__18113));
    InMux I__3981 (
            .O(N__18113),
            .I(N__18109));
    InMux I__3980 (
            .O(N__18112),
            .I(N__18106));
    LocalMux I__3979 (
            .O(N__18109),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__3978 (
            .O(N__18106),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__3977 (
            .O(N__18101),
            .I(N__18098));
    LocalMux I__3976 (
            .O(N__18098),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__3975 (
            .O(N__18095),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__3974 (
            .O(N__18092),
            .I(N__18088));
    InMux I__3973 (
            .O(N__18091),
            .I(N__18085));
    LocalMux I__3972 (
            .O(N__18088),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__3971 (
            .O(N__18085),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__3970 (
            .O(N__18080),
            .I(N__18077));
    InMux I__3969 (
            .O(N__18077),
            .I(N__18074));
    LocalMux I__3968 (
            .O(N__18074),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__3967 (
            .O(N__18071),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    CascadeMux I__3966 (
            .O(N__18068),
            .I(N__18065));
    InMux I__3965 (
            .O(N__18065),
            .I(N__18061));
    InMux I__3964 (
            .O(N__18064),
            .I(N__18058));
    LocalMux I__3963 (
            .O(N__18061),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__3962 (
            .O(N__18058),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__3961 (
            .O(N__18053),
            .I(N__18050));
    LocalMux I__3960 (
            .O(N__18050),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__3959 (
            .O(N__18047),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__3958 (
            .O(N__18044),
            .I(N__18041));
    LocalMux I__3957 (
            .O(N__18041),
            .I(N__18035));
    InMux I__3956 (
            .O(N__18040),
            .I(N__18032));
    CascadeMux I__3955 (
            .O(N__18039),
            .I(N__18028));
    CascadeMux I__3954 (
            .O(N__18038),
            .I(N__18025));
    Span4Mux_h I__3953 (
            .O(N__18035),
            .I(N__18019));
    LocalMux I__3952 (
            .O(N__18032),
            .I(N__18019));
    InMux I__3951 (
            .O(N__18031),
            .I(N__18016));
    InMux I__3950 (
            .O(N__18028),
            .I(N__18009));
    InMux I__3949 (
            .O(N__18025),
            .I(N__18009));
    InMux I__3948 (
            .O(N__18024),
            .I(N__18009));
    Span4Mux_h I__3947 (
            .O(N__18019),
            .I(N__18006));
    LocalMux I__3946 (
            .O(N__18016),
            .I(N__18001));
    LocalMux I__3945 (
            .O(N__18009),
            .I(N__18001));
    Odrv4 I__3944 (
            .O(N__18006),
            .I(\delay_measurement_inst.elapsed_time_hc_15 ));
    Odrv4 I__3943 (
            .O(N__18001),
            .I(\delay_measurement_inst.elapsed_time_hc_15 ));
    CascadeMux I__3942 (
            .O(N__17996),
            .I(N__17992));
    CascadeMux I__3941 (
            .O(N__17995),
            .I(N__17989));
    InMux I__3940 (
            .O(N__17992),
            .I(N__17986));
    InMux I__3939 (
            .O(N__17989),
            .I(N__17983));
    LocalMux I__3938 (
            .O(N__17986),
            .I(\delay_measurement_inst.N_84 ));
    LocalMux I__3937 (
            .O(N__17983),
            .I(\delay_measurement_inst.N_84 ));
    InMux I__3936 (
            .O(N__17978),
            .I(N__17975));
    LocalMux I__3935 (
            .O(N__17975),
            .I(N__17969));
    InMux I__3934 (
            .O(N__17974),
            .I(N__17966));
    InMux I__3933 (
            .O(N__17973),
            .I(N__17955));
    InMux I__3932 (
            .O(N__17972),
            .I(N__17955));
    Span4Mux_v I__3931 (
            .O(N__17969),
            .I(N__17950));
    LocalMux I__3930 (
            .O(N__17966),
            .I(N__17950));
    InMux I__3929 (
            .O(N__17965),
            .I(N__17945));
    InMux I__3928 (
            .O(N__17964),
            .I(N__17945));
    InMux I__3927 (
            .O(N__17963),
            .I(N__17936));
    InMux I__3926 (
            .O(N__17962),
            .I(N__17936));
    InMux I__3925 (
            .O(N__17961),
            .I(N__17936));
    InMux I__3924 (
            .O(N__17960),
            .I(N__17936));
    LocalMux I__3923 (
            .O(N__17955),
            .I(N__17933));
    Span4Mux_h I__3922 (
            .O(N__17950),
            .I(N__17926));
    LocalMux I__3921 (
            .O(N__17945),
            .I(N__17926));
    LocalMux I__3920 (
            .O(N__17936),
            .I(N__17926));
    Odrv4 I__3919 (
            .O(N__17933),
            .I(\delay_measurement_inst.N_40 ));
    Odrv4 I__3918 (
            .O(N__17926),
            .I(\delay_measurement_inst.N_40 ));
    CascadeMux I__3917 (
            .O(N__17921),
            .I(N__17917));
    InMux I__3916 (
            .O(N__17920),
            .I(N__17908));
    InMux I__3915 (
            .O(N__17917),
            .I(N__17908));
    InMux I__3914 (
            .O(N__17916),
            .I(N__17905));
    InMux I__3913 (
            .O(N__17915),
            .I(N__17902));
    InMux I__3912 (
            .O(N__17914),
            .I(N__17897));
    InMux I__3911 (
            .O(N__17913),
            .I(N__17897));
    LocalMux I__3910 (
            .O(N__17908),
            .I(N__17894));
    LocalMux I__3909 (
            .O(N__17905),
            .I(N__17891));
    LocalMux I__3908 (
            .O(N__17902),
            .I(N__17884));
    LocalMux I__3907 (
            .O(N__17897),
            .I(N__17884));
    Span4Mux_v I__3906 (
            .O(N__17894),
            .I(N__17884));
    Span4Mux_h I__3905 (
            .O(N__17891),
            .I(N__17881));
    Span4Mux_v I__3904 (
            .O(N__17884),
            .I(N__17875));
    Span4Mux_v I__3903 (
            .O(N__17881),
            .I(N__17872));
    InMux I__3902 (
            .O(N__17880),
            .I(N__17865));
    InMux I__3901 (
            .O(N__17879),
            .I(N__17865));
    InMux I__3900 (
            .O(N__17878),
            .I(N__17865));
    Odrv4 I__3899 (
            .O(N__17875),
            .I(measured_delay_hc_15));
    Odrv4 I__3898 (
            .O(N__17872),
            .I(measured_delay_hc_15));
    LocalMux I__3897 (
            .O(N__17865),
            .I(measured_delay_hc_15));
    InMux I__3896 (
            .O(N__17858),
            .I(N__17855));
    LocalMux I__3895 (
            .O(N__17855),
            .I(N__17851));
    InMux I__3894 (
            .O(N__17854),
            .I(N__17848));
    Span4Mux_h I__3893 (
            .O(N__17851),
            .I(N__17845));
    LocalMux I__3892 (
            .O(N__17848),
            .I(N__17842));
    Odrv4 I__3891 (
            .O(N__17845),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    Odrv4 I__3890 (
            .O(N__17842),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    CascadeMux I__3889 (
            .O(N__17837),
            .I(N__17834));
    InMux I__3888 (
            .O(N__17834),
            .I(N__17827));
    InMux I__3887 (
            .O(N__17833),
            .I(N__17827));
    CascadeMux I__3886 (
            .O(N__17832),
            .I(N__17822));
    LocalMux I__3885 (
            .O(N__17827),
            .I(N__17815));
    InMux I__3884 (
            .O(N__17826),
            .I(N__17806));
    InMux I__3883 (
            .O(N__17825),
            .I(N__17806));
    InMux I__3882 (
            .O(N__17822),
            .I(N__17806));
    InMux I__3881 (
            .O(N__17821),
            .I(N__17806));
    InMux I__3880 (
            .O(N__17820),
            .I(N__17799));
    InMux I__3879 (
            .O(N__17819),
            .I(N__17799));
    InMux I__3878 (
            .O(N__17818),
            .I(N__17799));
    Span4Mux_v I__3877 (
            .O(N__17815),
            .I(N__17789));
    LocalMux I__3876 (
            .O(N__17806),
            .I(N__17789));
    LocalMux I__3875 (
            .O(N__17799),
            .I(N__17786));
    InMux I__3874 (
            .O(N__17798),
            .I(N__17783));
    InMux I__3873 (
            .O(N__17797),
            .I(N__17780));
    InMux I__3872 (
            .O(N__17796),
            .I(N__17775));
    InMux I__3871 (
            .O(N__17795),
            .I(N__17775));
    InMux I__3870 (
            .O(N__17794),
            .I(N__17772));
    Span4Mux_v I__3869 (
            .O(N__17789),
            .I(N__17769));
    Span4Mux_h I__3868 (
            .O(N__17786),
            .I(N__17762));
    LocalMux I__3867 (
            .O(N__17783),
            .I(N__17762));
    LocalMux I__3866 (
            .O(N__17780),
            .I(N__17762));
    LocalMux I__3865 (
            .O(N__17775),
            .I(N__17759));
    LocalMux I__3864 (
            .O(N__17772),
            .I(N__17756));
    Span4Mux_h I__3863 (
            .O(N__17769),
            .I(N__17753));
    Span4Mux_h I__3862 (
            .O(N__17762),
            .I(N__17750));
    Span4Mux_v I__3861 (
            .O(N__17759),
            .I(N__17745));
    Span4Mux_v I__3860 (
            .O(N__17756),
            .I(N__17745));
    Odrv4 I__3859 (
            .O(N__17753),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    Odrv4 I__3858 (
            .O(N__17750),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    Odrv4 I__3857 (
            .O(N__17745),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    InMux I__3856 (
            .O(N__17738),
            .I(N__17735));
    LocalMux I__3855 (
            .O(N__17735),
            .I(N__17731));
    InMux I__3854 (
            .O(N__17734),
            .I(N__17728));
    Span4Mux_h I__3853 (
            .O(N__17731),
            .I(N__17725));
    LocalMux I__3852 (
            .O(N__17728),
            .I(N__17722));
    Odrv4 I__3851 (
            .O(N__17725),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    Odrv4 I__3850 (
            .O(N__17722),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__3849 (
            .O(N__17717),
            .I(N__17711));
    InMux I__3848 (
            .O(N__17716),
            .I(N__17711));
    LocalMux I__3847 (
            .O(N__17711),
            .I(N__17705));
    InMux I__3846 (
            .O(N__17710),
            .I(N__17702));
    InMux I__3845 (
            .O(N__17709),
            .I(N__17697));
    InMux I__3844 (
            .O(N__17708),
            .I(N__17697));
    Odrv4 I__3843 (
            .O(N__17705),
            .I(\delay_measurement_inst.N_48 ));
    LocalMux I__3842 (
            .O(N__17702),
            .I(\delay_measurement_inst.N_48 ));
    LocalMux I__3841 (
            .O(N__17697),
            .I(\delay_measurement_inst.N_48 ));
    CEMux I__3840 (
            .O(N__17690),
            .I(N__17687));
    LocalMux I__3839 (
            .O(N__17687),
            .I(N__17683));
    CEMux I__3838 (
            .O(N__17686),
            .I(N__17678));
    Span4Mux_h I__3837 (
            .O(N__17683),
            .I(N__17675));
    CEMux I__3836 (
            .O(N__17682),
            .I(N__17672));
    CEMux I__3835 (
            .O(N__17681),
            .I(N__17669));
    LocalMux I__3834 (
            .O(N__17678),
            .I(\delay_measurement_inst.N_54_i_0 ));
    Odrv4 I__3833 (
            .O(N__17675),
            .I(\delay_measurement_inst.N_54_i_0 ));
    LocalMux I__3832 (
            .O(N__17672),
            .I(\delay_measurement_inst.N_54_i_0 ));
    LocalMux I__3831 (
            .O(N__17669),
            .I(\delay_measurement_inst.N_54_i_0 ));
    SRMux I__3830 (
            .O(N__17660),
            .I(N__17645));
    SRMux I__3829 (
            .O(N__17659),
            .I(N__17645));
    SRMux I__3828 (
            .O(N__17658),
            .I(N__17645));
    SRMux I__3827 (
            .O(N__17657),
            .I(N__17645));
    SRMux I__3826 (
            .O(N__17656),
            .I(N__17645));
    GlobalMux I__3825 (
            .O(N__17645),
            .I(N__17642));
    gio2CtrlBuf I__3824 (
            .O(N__17642),
            .I(\delay_measurement_inst.N_32_g ));
    InMux I__3823 (
            .O(N__17639),
            .I(N__17627));
    InMux I__3822 (
            .O(N__17638),
            .I(N__17627));
    InMux I__3821 (
            .O(N__17637),
            .I(N__17627));
    InMux I__3820 (
            .O(N__17636),
            .I(N__17627));
    LocalMux I__3819 (
            .O(N__17627),
            .I(N__17614));
    InMux I__3818 (
            .O(N__17626),
            .I(N__17609));
    InMux I__3817 (
            .O(N__17625),
            .I(N__17609));
    InMux I__3816 (
            .O(N__17624),
            .I(N__17600));
    InMux I__3815 (
            .O(N__17623),
            .I(N__17600));
    InMux I__3814 (
            .O(N__17622),
            .I(N__17600));
    InMux I__3813 (
            .O(N__17621),
            .I(N__17600));
    InMux I__3812 (
            .O(N__17620),
            .I(N__17591));
    InMux I__3811 (
            .O(N__17619),
            .I(N__17591));
    InMux I__3810 (
            .O(N__17618),
            .I(N__17591));
    InMux I__3809 (
            .O(N__17617),
            .I(N__17591));
    Span4Mux_v I__3808 (
            .O(N__17614),
            .I(N__17578));
    LocalMux I__3807 (
            .O(N__17609),
            .I(N__17578));
    LocalMux I__3806 (
            .O(N__17600),
            .I(N__17578));
    LocalMux I__3805 (
            .O(N__17591),
            .I(N__17578));
    InMux I__3804 (
            .O(N__17590),
            .I(N__17561));
    InMux I__3803 (
            .O(N__17589),
            .I(N__17561));
    InMux I__3802 (
            .O(N__17588),
            .I(N__17561));
    InMux I__3801 (
            .O(N__17587),
            .I(N__17561));
    Span4Mux_v I__3800 (
            .O(N__17578),
            .I(N__17558));
    InMux I__3799 (
            .O(N__17577),
            .I(N__17549));
    InMux I__3798 (
            .O(N__17576),
            .I(N__17549));
    InMux I__3797 (
            .O(N__17575),
            .I(N__17549));
    InMux I__3796 (
            .O(N__17574),
            .I(N__17549));
    InMux I__3795 (
            .O(N__17573),
            .I(N__17540));
    InMux I__3794 (
            .O(N__17572),
            .I(N__17540));
    InMux I__3793 (
            .O(N__17571),
            .I(N__17540));
    InMux I__3792 (
            .O(N__17570),
            .I(N__17540));
    LocalMux I__3791 (
            .O(N__17561),
            .I(N__17533));
    Span4Mux_h I__3790 (
            .O(N__17558),
            .I(N__17526));
    LocalMux I__3789 (
            .O(N__17549),
            .I(N__17526));
    LocalMux I__3788 (
            .O(N__17540),
            .I(N__17526));
    InMux I__3787 (
            .O(N__17539),
            .I(N__17517));
    InMux I__3786 (
            .O(N__17538),
            .I(N__17517));
    InMux I__3785 (
            .O(N__17537),
            .I(N__17517));
    InMux I__3784 (
            .O(N__17536),
            .I(N__17517));
    Span4Mux_v I__3783 (
            .O(N__17533),
            .I(N__17512));
    Span4Mux_h I__3782 (
            .O(N__17526),
            .I(N__17512));
    LocalMux I__3781 (
            .O(N__17517),
            .I(N__17509));
    Span4Mux_h I__3780 (
            .O(N__17512),
            .I(N__17506));
    Odrv12 I__3779 (
            .O(N__17509),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__3778 (
            .O(N__17506),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    CEMux I__3777 (
            .O(N__17501),
            .I(N__17495));
    CEMux I__3776 (
            .O(N__17500),
            .I(N__17492));
    CEMux I__3775 (
            .O(N__17499),
            .I(N__17489));
    CEMux I__3774 (
            .O(N__17498),
            .I(N__17486));
    LocalMux I__3773 (
            .O(N__17495),
            .I(N__17481));
    LocalMux I__3772 (
            .O(N__17492),
            .I(N__17481));
    LocalMux I__3771 (
            .O(N__17489),
            .I(N__17478));
    LocalMux I__3770 (
            .O(N__17486),
            .I(N__17475));
    Span4Mux_v I__3769 (
            .O(N__17481),
            .I(N__17472));
    Span4Mux_h I__3768 (
            .O(N__17478),
            .I(N__17469));
    Sp12to4 I__3767 (
            .O(N__17475),
            .I(N__17466));
    Span4Mux_h I__3766 (
            .O(N__17472),
            .I(N__17463));
    Span4Mux_h I__3765 (
            .O(N__17469),
            .I(N__17460));
    Odrv12 I__3764 (
            .O(N__17466),
            .I(\delay_measurement_inst.delay_hc_timer.N_179_i_g ));
    Odrv4 I__3763 (
            .O(N__17463),
            .I(\delay_measurement_inst.delay_hc_timer.N_179_i_g ));
    Odrv4 I__3762 (
            .O(N__17460),
            .I(\delay_measurement_inst.delay_hc_timer.N_179_i_g ));
    InMux I__3761 (
            .O(N__17453),
            .I(N__17448));
    InMux I__3760 (
            .O(N__17452),
            .I(N__17445));
    InMux I__3759 (
            .O(N__17451),
            .I(N__17442));
    LocalMux I__3758 (
            .O(N__17448),
            .I(N__17439));
    LocalMux I__3757 (
            .O(N__17445),
            .I(N__17435));
    LocalMux I__3756 (
            .O(N__17442),
            .I(N__17432));
    Span4Mux_v I__3755 (
            .O(N__17439),
            .I(N__17429));
    InMux I__3754 (
            .O(N__17438),
            .I(N__17426));
    Span4Mux_h I__3753 (
            .O(N__17435),
            .I(N__17421));
    Span4Mux_v I__3752 (
            .O(N__17432),
            .I(N__17421));
    Odrv4 I__3751 (
            .O(N__17429),
            .I(measured_delay_hc_2));
    LocalMux I__3750 (
            .O(N__17426),
            .I(measured_delay_hc_2));
    Odrv4 I__3749 (
            .O(N__17421),
            .I(measured_delay_hc_2));
    InMux I__3748 (
            .O(N__17414),
            .I(N__17411));
    LocalMux I__3747 (
            .O(N__17411),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto6Z0Z_0 ));
    CascadeMux I__3746 (
            .O(N__17408),
            .I(N__17404));
    CascadeMux I__3745 (
            .O(N__17407),
            .I(N__17401));
    InMux I__3744 (
            .O(N__17404),
            .I(N__17396));
    InMux I__3743 (
            .O(N__17401),
            .I(N__17393));
    CascadeMux I__3742 (
            .O(N__17400),
            .I(N__17390));
    InMux I__3741 (
            .O(N__17399),
            .I(N__17387));
    LocalMux I__3740 (
            .O(N__17396),
            .I(N__17384));
    LocalMux I__3739 (
            .O(N__17393),
            .I(N__17381));
    InMux I__3738 (
            .O(N__17390),
            .I(N__17378));
    LocalMux I__3737 (
            .O(N__17387),
            .I(N__17375));
    Span4Mux_v I__3736 (
            .O(N__17384),
            .I(N__17370));
    Span4Mux_h I__3735 (
            .O(N__17381),
            .I(N__17370));
    LocalMux I__3734 (
            .O(N__17378),
            .I(measured_delay_hc_3));
    Odrv4 I__3733 (
            .O(N__17375),
            .I(measured_delay_hc_3));
    Odrv4 I__3732 (
            .O(N__17370),
            .I(measured_delay_hc_3));
    CascadeMux I__3731 (
            .O(N__17363),
            .I(N__17359));
    InMux I__3730 (
            .O(N__17362),
            .I(N__17356));
    InMux I__3729 (
            .O(N__17359),
            .I(N__17352));
    LocalMux I__3728 (
            .O(N__17356),
            .I(N__17349));
    InMux I__3727 (
            .O(N__17355),
            .I(N__17346));
    LocalMux I__3726 (
            .O(N__17352),
            .I(N__17342));
    Span4Mux_v I__3725 (
            .O(N__17349),
            .I(N__17337));
    LocalMux I__3724 (
            .O(N__17346),
            .I(N__17337));
    InMux I__3723 (
            .O(N__17345),
            .I(N__17334));
    Odrv4 I__3722 (
            .O(N__17342),
            .I(measured_delay_hc_4));
    Odrv4 I__3721 (
            .O(N__17337),
            .I(measured_delay_hc_4));
    LocalMux I__3720 (
            .O(N__17334),
            .I(measured_delay_hc_4));
    InMux I__3719 (
            .O(N__17327),
            .I(N__17324));
    LocalMux I__3718 (
            .O(N__17324),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_4 ));
    InMux I__3717 (
            .O(N__17321),
            .I(N__17317));
    InMux I__3716 (
            .O(N__17320),
            .I(N__17314));
    LocalMux I__3715 (
            .O(N__17317),
            .I(N__17310));
    LocalMux I__3714 (
            .O(N__17314),
            .I(N__17306));
    InMux I__3713 (
            .O(N__17313),
            .I(N__17303));
    Span12Mux_h I__3712 (
            .O(N__17310),
            .I(N__17300));
    InMux I__3711 (
            .O(N__17309),
            .I(N__17297));
    Span4Mux_v I__3710 (
            .O(N__17306),
            .I(N__17292));
    LocalMux I__3709 (
            .O(N__17303),
            .I(N__17292));
    Odrv12 I__3708 (
            .O(N__17300),
            .I(measured_delay_hc_12));
    LocalMux I__3707 (
            .O(N__17297),
            .I(measured_delay_hc_12));
    Odrv4 I__3706 (
            .O(N__17292),
            .I(measured_delay_hc_12));
    CascadeMux I__3705 (
            .O(N__17285),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt19_0_cascade_ ));
    InMux I__3704 (
            .O(N__17282),
            .I(N__17279));
    LocalMux I__3703 (
            .O(N__17279),
            .I(N__17275));
    InMux I__3702 (
            .O(N__17278),
            .I(N__17272));
    Span4Mux_h I__3701 (
            .O(N__17275),
            .I(N__17269));
    LocalMux I__3700 (
            .O(N__17272),
            .I(N__17266));
    Span4Mux_v I__3699 (
            .O(N__17269),
            .I(N__17261));
    Span4Mux_h I__3698 (
            .O(N__17266),
            .I(N__17258));
    InMux I__3697 (
            .O(N__17265),
            .I(N__17255));
    InMux I__3696 (
            .O(N__17264),
            .I(N__17252));
    Odrv4 I__3695 (
            .O(N__17261),
            .I(measured_delay_hc_11));
    Odrv4 I__3694 (
            .O(N__17258),
            .I(measured_delay_hc_11));
    LocalMux I__3693 (
            .O(N__17255),
            .I(measured_delay_hc_11));
    LocalMux I__3692 (
            .O(N__17252),
            .I(measured_delay_hc_11));
    CascadeMux I__3691 (
            .O(N__17243),
            .I(N__17239));
    CascadeMux I__3690 (
            .O(N__17242),
            .I(N__17235));
    InMux I__3689 (
            .O(N__17239),
            .I(N__17229));
    InMux I__3688 (
            .O(N__17238),
            .I(N__17229));
    InMux I__3687 (
            .O(N__17235),
            .I(N__17224));
    InMux I__3686 (
            .O(N__17234),
            .I(N__17224));
    LocalMux I__3685 (
            .O(N__17229),
            .I(N__17221));
    LocalMux I__3684 (
            .O(N__17224),
            .I(N__17218));
    Span4Mux_h I__3683 (
            .O(N__17221),
            .I(N__17214));
    Span4Mux_h I__3682 (
            .O(N__17218),
            .I(N__17211));
    InMux I__3681 (
            .O(N__17217),
            .I(N__17208));
    Odrv4 I__3680 (
            .O(N__17214),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9 ));
    Odrv4 I__3679 (
            .O(N__17211),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9 ));
    LocalMux I__3678 (
            .O(N__17208),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9 ));
    InMux I__3677 (
            .O(N__17201),
            .I(N__17198));
    LocalMux I__3676 (
            .O(N__17198),
            .I(N__17195));
    Span4Mux_v I__3675 (
            .O(N__17195),
            .I(N__17192));
    Span4Mux_h I__3674 (
            .O(N__17192),
            .I(N__17189));
    Odrv4 I__3673 (
            .O(N__17189),
            .I(il_max_comp1_D1));
    SRMux I__3672 (
            .O(N__17186),
            .I(N__17180));
    SRMux I__3671 (
            .O(N__17185),
            .I(N__17176));
    SRMux I__3670 (
            .O(N__17184),
            .I(N__17173));
    SRMux I__3669 (
            .O(N__17183),
            .I(N__17169));
    LocalMux I__3668 (
            .O(N__17180),
            .I(N__17166));
    SRMux I__3667 (
            .O(N__17179),
            .I(N__17163));
    LocalMux I__3666 (
            .O(N__17176),
            .I(N__17160));
    LocalMux I__3665 (
            .O(N__17173),
            .I(N__17157));
    SRMux I__3664 (
            .O(N__17172),
            .I(N__17154));
    LocalMux I__3663 (
            .O(N__17169),
            .I(N__17151));
    Span4Mux_v I__3662 (
            .O(N__17166),
            .I(N__17146));
    LocalMux I__3661 (
            .O(N__17163),
            .I(N__17146));
    Span4Mux_v I__3660 (
            .O(N__17160),
            .I(N__17142));
    Span4Mux_h I__3659 (
            .O(N__17157),
            .I(N__17137));
    LocalMux I__3658 (
            .O(N__17154),
            .I(N__17137));
    Span4Mux_h I__3657 (
            .O(N__17151),
            .I(N__17132));
    Span4Mux_h I__3656 (
            .O(N__17146),
            .I(N__17132));
    InMux I__3655 (
            .O(N__17145),
            .I(N__17129));
    Odrv4 I__3654 (
            .O(N__17142),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31 ));
    Odrv4 I__3653 (
            .O(N__17137),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31 ));
    Odrv4 I__3652 (
            .O(N__17132),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31 ));
    LocalMux I__3651 (
            .O(N__17129),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31 ));
    InMux I__3650 (
            .O(N__17120),
            .I(N__17117));
    LocalMux I__3649 (
            .O(N__17117),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_7_9 ));
    InMux I__3648 (
            .O(N__17114),
            .I(N__17111));
    LocalMux I__3647 (
            .O(N__17111),
            .I(\delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_4 ));
    InMux I__3646 (
            .O(N__17108),
            .I(N__17105));
    LocalMux I__3645 (
            .O(N__17105),
            .I(N__17100));
    InMux I__3644 (
            .O(N__17104),
            .I(N__17095));
    InMux I__3643 (
            .O(N__17103),
            .I(N__17095));
    Odrv4 I__3642 (
            .O(N__17100),
            .I(\delay_measurement_inst.delay_tr_timer.N_127 ));
    LocalMux I__3641 (
            .O(N__17095),
            .I(\delay_measurement_inst.delay_tr_timer.N_127 ));
    InMux I__3640 (
            .O(N__17090),
            .I(N__17087));
    LocalMux I__3639 (
            .O(N__17087),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_6_9 ));
    InMux I__3638 (
            .O(N__17084),
            .I(N__17081));
    LocalMux I__3637 (
            .O(N__17081),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_0_9 ));
    InMux I__3636 (
            .O(N__17078),
            .I(N__17075));
    LocalMux I__3635 (
            .O(N__17075),
            .I(N__17072));
    Glb2LocalMux I__3634 (
            .O(N__17072),
            .I(N__17069));
    GlobalMux I__3633 (
            .O(N__17069),
            .I(clk_12mhz));
    IoInMux I__3632 (
            .O(N__17066),
            .I(N__17063));
    LocalMux I__3631 (
            .O(N__17063),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__3630 (
            .O(N__17060),
            .I(N__17057));
    LocalMux I__3629 (
            .O(N__17057),
            .I(delay_hc_d2));
    InMux I__3628 (
            .O(N__17054),
            .I(N__17051));
    LocalMux I__3627 (
            .O(N__17051),
            .I(\delay_measurement_inst.hc_syncZ0Z_0 ));
    InMux I__3626 (
            .O(N__17048),
            .I(N__17045));
    LocalMux I__3625 (
            .O(N__17045),
            .I(N__17041));
    InMux I__3624 (
            .O(N__17044),
            .I(N__17036));
    Span4Mux_h I__3623 (
            .O(N__17041),
            .I(N__17033));
    InMux I__3622 (
            .O(N__17040),
            .I(N__17030));
    InMux I__3621 (
            .O(N__17039),
            .I(N__17027));
    LocalMux I__3620 (
            .O(N__17036),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__3619 (
            .O(N__17033),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__3618 (
            .O(N__17030),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__3617 (
            .O(N__17027),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    CascadeMux I__3616 (
            .O(N__17018),
            .I(N__17015));
    InMux I__3615 (
            .O(N__17015),
            .I(N__17012));
    LocalMux I__3614 (
            .O(N__17012),
            .I(N__17009));
    Span4Mux_h I__3613 (
            .O(N__17009),
            .I(N__17006));
    Span4Mux_h I__3612 (
            .O(N__17006),
            .I(N__17003));
    Odrv4 I__3611 (
            .O(N__17003),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    InMux I__3610 (
            .O(N__17000),
            .I(N__16996));
    InMux I__3609 (
            .O(N__16999),
            .I(N__16993));
    LocalMux I__3608 (
            .O(N__16996),
            .I(N__16990));
    LocalMux I__3607 (
            .O(N__16993),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    Odrv4 I__3606 (
            .O(N__16990),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    InMux I__3605 (
            .O(N__16985),
            .I(N__16977));
    InMux I__3604 (
            .O(N__16984),
            .I(N__16971));
    InMux I__3603 (
            .O(N__16983),
            .I(N__16968));
    InMux I__3602 (
            .O(N__16982),
            .I(N__16961));
    InMux I__3601 (
            .O(N__16981),
            .I(N__16961));
    InMux I__3600 (
            .O(N__16980),
            .I(N__16961));
    LocalMux I__3599 (
            .O(N__16977),
            .I(N__16958));
    InMux I__3598 (
            .O(N__16976),
            .I(N__16955));
    InMux I__3597 (
            .O(N__16975),
            .I(N__16952));
    InMux I__3596 (
            .O(N__16974),
            .I(N__16949));
    LocalMux I__3595 (
            .O(N__16971),
            .I(\delay_measurement_inst.N_201 ));
    LocalMux I__3594 (
            .O(N__16968),
            .I(\delay_measurement_inst.N_201 ));
    LocalMux I__3593 (
            .O(N__16961),
            .I(\delay_measurement_inst.N_201 ));
    Odrv4 I__3592 (
            .O(N__16958),
            .I(\delay_measurement_inst.N_201 ));
    LocalMux I__3591 (
            .O(N__16955),
            .I(\delay_measurement_inst.N_201 ));
    LocalMux I__3590 (
            .O(N__16952),
            .I(\delay_measurement_inst.N_201 ));
    LocalMux I__3589 (
            .O(N__16949),
            .I(\delay_measurement_inst.N_201 ));
    InMux I__3588 (
            .O(N__16934),
            .I(N__16930));
    InMux I__3587 (
            .O(N__16933),
            .I(N__16927));
    LocalMux I__3586 (
            .O(N__16930),
            .I(N__16920));
    LocalMux I__3585 (
            .O(N__16927),
            .I(N__16920));
    InMux I__3584 (
            .O(N__16926),
            .I(N__16917));
    InMux I__3583 (
            .O(N__16925),
            .I(N__16914));
    Span4Mux_v I__3582 (
            .O(N__16920),
            .I(N__16911));
    LocalMux I__3581 (
            .O(N__16917),
            .I(N__16908));
    LocalMux I__3580 (
            .O(N__16914),
            .I(N__16905));
    Span4Mux_h I__3579 (
            .O(N__16911),
            .I(N__16900));
    Span4Mux_v I__3578 (
            .O(N__16908),
            .I(N__16900));
    Span4Mux_h I__3577 (
            .O(N__16905),
            .I(N__16897));
    Odrv4 I__3576 (
            .O(N__16900),
            .I(measured_delay_tr_19));
    Odrv4 I__3575 (
            .O(N__16897),
            .I(measured_delay_tr_19));
    CEMux I__3574 (
            .O(N__16892),
            .I(N__16888));
    CEMux I__3573 (
            .O(N__16891),
            .I(N__16883));
    LocalMux I__3572 (
            .O(N__16888),
            .I(N__16880));
    CEMux I__3571 (
            .O(N__16887),
            .I(N__16877));
    CEMux I__3570 (
            .O(N__16886),
            .I(N__16874));
    LocalMux I__3569 (
            .O(N__16883),
            .I(N__16871));
    Span4Mux_h I__3568 (
            .O(N__16880),
            .I(N__16866));
    LocalMux I__3567 (
            .O(N__16877),
            .I(N__16866));
    LocalMux I__3566 (
            .O(N__16874),
            .I(N__16863));
    Span4Mux_h I__3565 (
            .O(N__16871),
            .I(N__16860));
    Span4Mux_h I__3564 (
            .O(N__16866),
            .I(N__16855));
    Span4Mux_h I__3563 (
            .O(N__16863),
            .I(N__16855));
    Odrv4 I__3562 (
            .O(N__16860),
            .I(\delay_measurement_inst.N_134_i_0 ));
    Odrv4 I__3561 (
            .O(N__16855),
            .I(\delay_measurement_inst.N_134_i_0 ));
    CascadeMux I__3560 (
            .O(N__16850),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ));
    InMux I__3559 (
            .O(N__16847),
            .I(N__16843));
    InMux I__3558 (
            .O(N__16846),
            .I(N__16840));
    LocalMux I__3557 (
            .O(N__16843),
            .I(N__16837));
    LocalMux I__3556 (
            .O(N__16840),
            .I(N__16832));
    Span4Mux_h I__3555 (
            .O(N__16837),
            .I(N__16829));
    InMux I__3554 (
            .O(N__16836),
            .I(N__16826));
    InMux I__3553 (
            .O(N__16835),
            .I(N__16823));
    Odrv4 I__3552 (
            .O(N__16832),
            .I(measured_delay_hc_6));
    Odrv4 I__3551 (
            .O(N__16829),
            .I(measured_delay_hc_6));
    LocalMux I__3550 (
            .O(N__16826),
            .I(measured_delay_hc_6));
    LocalMux I__3549 (
            .O(N__16823),
            .I(measured_delay_hc_6));
    InMux I__3548 (
            .O(N__16814),
            .I(N__16811));
    LocalMux I__3547 (
            .O(N__16811),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ));
    InMux I__3546 (
            .O(N__16808),
            .I(N__16805));
    LocalMux I__3545 (
            .O(N__16805),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__3544 (
            .O(N__16802),
            .I(N__16798));
    InMux I__3543 (
            .O(N__16801),
            .I(N__16795));
    LocalMux I__3542 (
            .O(N__16798),
            .I(N__16792));
    LocalMux I__3541 (
            .O(N__16795),
            .I(N__16786));
    Span4Mux_v I__3540 (
            .O(N__16792),
            .I(N__16783));
    InMux I__3539 (
            .O(N__16791),
            .I(N__16776));
    InMux I__3538 (
            .O(N__16790),
            .I(N__16776));
    InMux I__3537 (
            .O(N__16789),
            .I(N__16776));
    Odrv12 I__3536 (
            .O(N__16786),
            .I(measured_delay_hc_9));
    Odrv4 I__3535 (
            .O(N__16783),
            .I(measured_delay_hc_9));
    LocalMux I__3534 (
            .O(N__16776),
            .I(measured_delay_hc_9));
    InMux I__3533 (
            .O(N__16769),
            .I(N__16766));
    LocalMux I__3532 (
            .O(N__16766),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__3531 (
            .O(N__16763),
            .I(N__16760));
    LocalMux I__3530 (
            .O(N__16760),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__3529 (
            .O(N__16757),
            .I(N__16753));
    CascadeMux I__3528 (
            .O(N__16756),
            .I(N__16750));
    InMux I__3527 (
            .O(N__16753),
            .I(N__16747));
    InMux I__3526 (
            .O(N__16750),
            .I(N__16744));
    LocalMux I__3525 (
            .O(N__16747),
            .I(N__16740));
    LocalMux I__3524 (
            .O(N__16744),
            .I(N__16737));
    InMux I__3523 (
            .O(N__16743),
            .I(N__16734));
    Odrv4 I__3522 (
            .O(N__16740),
            .I(measured_delay_hc_13));
    Odrv12 I__3521 (
            .O(N__16737),
            .I(measured_delay_hc_13));
    LocalMux I__3520 (
            .O(N__16734),
            .I(measured_delay_hc_13));
    InMux I__3519 (
            .O(N__16727),
            .I(N__16724));
    LocalMux I__3518 (
            .O(N__16724),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__3517 (
            .O(N__16721),
            .I(N__16700));
    InMux I__3516 (
            .O(N__16720),
            .I(N__16700));
    InMux I__3515 (
            .O(N__16719),
            .I(N__16700));
    InMux I__3514 (
            .O(N__16718),
            .I(N__16700));
    InMux I__3513 (
            .O(N__16717),
            .I(N__16700));
    InMux I__3512 (
            .O(N__16716),
            .I(N__16697));
    InMux I__3511 (
            .O(N__16715),
            .I(N__16686));
    InMux I__3510 (
            .O(N__16714),
            .I(N__16686));
    InMux I__3509 (
            .O(N__16713),
            .I(N__16686));
    InMux I__3508 (
            .O(N__16712),
            .I(N__16686));
    InMux I__3507 (
            .O(N__16711),
            .I(N__16686));
    LocalMux I__3506 (
            .O(N__16700),
            .I(N__16672));
    LocalMux I__3505 (
            .O(N__16697),
            .I(N__16667));
    LocalMux I__3504 (
            .O(N__16686),
            .I(N__16667));
    InMux I__3503 (
            .O(N__16685),
            .I(N__16656));
    InMux I__3502 (
            .O(N__16684),
            .I(N__16656));
    InMux I__3501 (
            .O(N__16683),
            .I(N__16656));
    InMux I__3500 (
            .O(N__16682),
            .I(N__16656));
    InMux I__3499 (
            .O(N__16681),
            .I(N__16656));
    InMux I__3498 (
            .O(N__16680),
            .I(N__16643));
    InMux I__3497 (
            .O(N__16679),
            .I(N__16643));
    InMux I__3496 (
            .O(N__16678),
            .I(N__16643));
    InMux I__3495 (
            .O(N__16677),
            .I(N__16643));
    InMux I__3494 (
            .O(N__16676),
            .I(N__16643));
    InMux I__3493 (
            .O(N__16675),
            .I(N__16643));
    Span4Mux_v I__3492 (
            .O(N__16672),
            .I(N__16639));
    Span4Mux_v I__3491 (
            .O(N__16667),
            .I(N__16632));
    LocalMux I__3490 (
            .O(N__16656),
            .I(N__16632));
    LocalMux I__3489 (
            .O(N__16643),
            .I(N__16632));
    InMux I__3488 (
            .O(N__16642),
            .I(N__16629));
    Odrv4 I__3487 (
            .O(N__16639),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt15 ));
    Odrv4 I__3486 (
            .O(N__16632),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt15 ));
    LocalMux I__3485 (
            .O(N__16629),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt15 ));
    CascadeMux I__3484 (
            .O(N__16622),
            .I(N__16617));
    CascadeMux I__3483 (
            .O(N__16621),
            .I(N__16614));
    CascadeMux I__3482 (
            .O(N__16620),
            .I(N__16611));
    InMux I__3481 (
            .O(N__16617),
            .I(N__16590));
    InMux I__3480 (
            .O(N__16614),
            .I(N__16590));
    InMux I__3479 (
            .O(N__16611),
            .I(N__16590));
    InMux I__3478 (
            .O(N__16610),
            .I(N__16590));
    InMux I__3477 (
            .O(N__16609),
            .I(N__16590));
    CascadeMux I__3476 (
            .O(N__16608),
            .I(N__16587));
    CascadeMux I__3475 (
            .O(N__16607),
            .I(N__16584));
    CascadeMux I__3474 (
            .O(N__16606),
            .I(N__16581));
    InMux I__3473 (
            .O(N__16605),
            .I(N__16576));
    InMux I__3472 (
            .O(N__16604),
            .I(N__16567));
    InMux I__3471 (
            .O(N__16603),
            .I(N__16567));
    InMux I__3470 (
            .O(N__16602),
            .I(N__16567));
    InMux I__3469 (
            .O(N__16601),
            .I(N__16567));
    LocalMux I__3468 (
            .O(N__16590),
            .I(N__16559));
    InMux I__3467 (
            .O(N__16587),
            .I(N__16548));
    InMux I__3466 (
            .O(N__16584),
            .I(N__16548));
    InMux I__3465 (
            .O(N__16581),
            .I(N__16548));
    InMux I__3464 (
            .O(N__16580),
            .I(N__16548));
    InMux I__3463 (
            .O(N__16579),
            .I(N__16548));
    LocalMux I__3462 (
            .O(N__16576),
            .I(N__16545));
    LocalMux I__3461 (
            .O(N__16567),
            .I(N__16542));
    InMux I__3460 (
            .O(N__16566),
            .I(N__16531));
    InMux I__3459 (
            .O(N__16565),
            .I(N__16531));
    InMux I__3458 (
            .O(N__16564),
            .I(N__16531));
    InMux I__3457 (
            .O(N__16563),
            .I(N__16531));
    InMux I__3456 (
            .O(N__16562),
            .I(N__16531));
    Span4Mux_v I__3455 (
            .O(N__16559),
            .I(N__16528));
    LocalMux I__3454 (
            .O(N__16548),
            .I(N__16521));
    Span4Mux_v I__3453 (
            .O(N__16545),
            .I(N__16521));
    Span4Mux_v I__3452 (
            .O(N__16542),
            .I(N__16521));
    LocalMux I__3451 (
            .O(N__16531),
            .I(\phase_controller_inst1.stoper_hc.un3_start ));
    Odrv4 I__3450 (
            .O(N__16528),
            .I(\phase_controller_inst1.stoper_hc.un3_start ));
    Odrv4 I__3449 (
            .O(N__16521),
            .I(\phase_controller_inst1.stoper_hc.un3_start ));
    InMux I__3448 (
            .O(N__16514),
            .I(N__16510));
    InMux I__3447 (
            .O(N__16513),
            .I(N__16507));
    LocalMux I__3446 (
            .O(N__16510),
            .I(N__16503));
    LocalMux I__3445 (
            .O(N__16507),
            .I(N__16500));
    InMux I__3444 (
            .O(N__16506),
            .I(N__16497));
    Odrv12 I__3443 (
            .O(N__16503),
            .I(measured_delay_hc_10));
    Odrv4 I__3442 (
            .O(N__16500),
            .I(measured_delay_hc_10));
    LocalMux I__3441 (
            .O(N__16497),
            .I(measured_delay_hc_10));
    InMux I__3440 (
            .O(N__16490),
            .I(N__16487));
    LocalMux I__3439 (
            .O(N__16487),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__3438 (
            .O(N__16484),
            .I(N__16481));
    LocalMux I__3437 (
            .O(N__16481),
            .I(N__16477));
    InMux I__3436 (
            .O(N__16480),
            .I(N__16474));
    Span4Mux_v I__3435 (
            .O(N__16477),
            .I(N__16469));
    LocalMux I__3434 (
            .O(N__16474),
            .I(N__16469));
    Span4Mux_v I__3433 (
            .O(N__16469),
            .I(N__16464));
    InMux I__3432 (
            .O(N__16468),
            .I(N__16461));
    InMux I__3431 (
            .O(N__16467),
            .I(N__16458));
    Odrv4 I__3430 (
            .O(N__16464),
            .I(measured_delay_hc_14));
    LocalMux I__3429 (
            .O(N__16461),
            .I(measured_delay_hc_14));
    LocalMux I__3428 (
            .O(N__16458),
            .I(measured_delay_hc_14));
    InMux I__3427 (
            .O(N__16451),
            .I(N__16448));
    LocalMux I__3426 (
            .O(N__16448),
            .I(N__16445));
    Odrv4 I__3425 (
            .O(N__16445),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__3424 (
            .O(N__16442),
            .I(N__16431));
    CascadeMux I__3423 (
            .O(N__16441),
            .I(N__16425));
    CascadeMux I__3422 (
            .O(N__16440),
            .I(N__16422));
    CascadeMux I__3421 (
            .O(N__16439),
            .I(N__16419));
    CascadeMux I__3420 (
            .O(N__16438),
            .I(N__16416));
    InMux I__3419 (
            .O(N__16437),
            .I(N__16401));
    InMux I__3418 (
            .O(N__16436),
            .I(N__16401));
    InMux I__3417 (
            .O(N__16435),
            .I(N__16401));
    InMux I__3416 (
            .O(N__16434),
            .I(N__16401));
    InMux I__3415 (
            .O(N__16431),
            .I(N__16401));
    InMux I__3414 (
            .O(N__16430),
            .I(N__16393));
    InMux I__3413 (
            .O(N__16429),
            .I(N__16393));
    InMux I__3412 (
            .O(N__16428),
            .I(N__16380));
    InMux I__3411 (
            .O(N__16425),
            .I(N__16380));
    InMux I__3410 (
            .O(N__16422),
            .I(N__16380));
    InMux I__3409 (
            .O(N__16419),
            .I(N__16380));
    InMux I__3408 (
            .O(N__16416),
            .I(N__16380));
    InMux I__3407 (
            .O(N__16415),
            .I(N__16380));
    CascadeMux I__3406 (
            .O(N__16414),
            .I(N__16377));
    CascadeMux I__3405 (
            .O(N__16413),
            .I(N__16374));
    CascadeMux I__3404 (
            .O(N__16412),
            .I(N__16367));
    LocalMux I__3403 (
            .O(N__16401),
            .I(N__16363));
    CascadeMux I__3402 (
            .O(N__16400),
            .I(N__16360));
    CascadeMux I__3401 (
            .O(N__16399),
            .I(N__16357));
    CascadeMux I__3400 (
            .O(N__16398),
            .I(N__16352));
    LocalMux I__3399 (
            .O(N__16393),
            .I(N__16347));
    LocalMux I__3398 (
            .O(N__16380),
            .I(N__16347));
    InMux I__3397 (
            .O(N__16377),
            .I(N__16330));
    InMux I__3396 (
            .O(N__16374),
            .I(N__16330));
    InMux I__3395 (
            .O(N__16373),
            .I(N__16330));
    InMux I__3394 (
            .O(N__16372),
            .I(N__16330));
    InMux I__3393 (
            .O(N__16371),
            .I(N__16330));
    InMux I__3392 (
            .O(N__16370),
            .I(N__16330));
    InMux I__3391 (
            .O(N__16367),
            .I(N__16330));
    InMux I__3390 (
            .O(N__16366),
            .I(N__16330));
    Span4Mux_h I__3389 (
            .O(N__16363),
            .I(N__16326));
    InMux I__3388 (
            .O(N__16360),
            .I(N__16315));
    InMux I__3387 (
            .O(N__16357),
            .I(N__16315));
    InMux I__3386 (
            .O(N__16356),
            .I(N__16315));
    InMux I__3385 (
            .O(N__16355),
            .I(N__16315));
    InMux I__3384 (
            .O(N__16352),
            .I(N__16315));
    Span4Mux_v I__3383 (
            .O(N__16347),
            .I(N__16310));
    LocalMux I__3382 (
            .O(N__16330),
            .I(N__16310));
    InMux I__3381 (
            .O(N__16329),
            .I(N__16307));
    Odrv4 I__3380 (
            .O(N__16326),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    LocalMux I__3379 (
            .O(N__16315),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    Odrv4 I__3378 (
            .O(N__16310),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    LocalMux I__3377 (
            .O(N__16307),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    InMux I__3376 (
            .O(N__16298),
            .I(N__16295));
    LocalMux I__3375 (
            .O(N__16295),
            .I(N__16292));
    Odrv4 I__3374 (
            .O(N__16292),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__3373 (
            .O(N__16289),
            .I(N__16286));
    LocalMux I__3372 (
            .O(N__16286),
            .I(N__16280));
    InMux I__3371 (
            .O(N__16285),
            .I(N__16277));
    InMux I__3370 (
            .O(N__16284),
            .I(N__16272));
    InMux I__3369 (
            .O(N__16283),
            .I(N__16272));
    Odrv4 I__3368 (
            .O(N__16280),
            .I(measured_delay_hc_5));
    LocalMux I__3367 (
            .O(N__16277),
            .I(measured_delay_hc_5));
    LocalMux I__3366 (
            .O(N__16272),
            .I(measured_delay_hc_5));
    InMux I__3365 (
            .O(N__16265),
            .I(N__16262));
    LocalMux I__3364 (
            .O(N__16262),
            .I(N__16256));
    InMux I__3363 (
            .O(N__16261),
            .I(N__16253));
    InMux I__3362 (
            .O(N__16260),
            .I(N__16248));
    InMux I__3361 (
            .O(N__16259),
            .I(N__16248));
    Span4Mux_v I__3360 (
            .O(N__16256),
            .I(N__16245));
    LocalMux I__3359 (
            .O(N__16253),
            .I(N__16242));
    LocalMux I__3358 (
            .O(N__16248),
            .I(N__16239));
    Odrv4 I__3357 (
            .O(N__16245),
            .I(measured_delay_hc_16));
    Odrv4 I__3356 (
            .O(N__16242),
            .I(measured_delay_hc_16));
    Odrv4 I__3355 (
            .O(N__16239),
            .I(measured_delay_hc_16));
    InMux I__3354 (
            .O(N__16232),
            .I(N__16229));
    LocalMux I__3353 (
            .O(N__16229),
            .I(N__16223));
    InMux I__3352 (
            .O(N__16228),
            .I(N__16220));
    InMux I__3351 (
            .O(N__16227),
            .I(N__16215));
    InMux I__3350 (
            .O(N__16226),
            .I(N__16215));
    Span4Mux_v I__3349 (
            .O(N__16223),
            .I(N__16212));
    LocalMux I__3348 (
            .O(N__16220),
            .I(N__16209));
    LocalMux I__3347 (
            .O(N__16215),
            .I(N__16206));
    Odrv4 I__3346 (
            .O(N__16212),
            .I(measured_delay_hc_19));
    Odrv4 I__3345 (
            .O(N__16209),
            .I(measured_delay_hc_19));
    Odrv4 I__3344 (
            .O(N__16206),
            .I(measured_delay_hc_19));
    InMux I__3343 (
            .O(N__16199),
            .I(N__16196));
    LocalMux I__3342 (
            .O(N__16196),
            .I(N__16190));
    InMux I__3341 (
            .O(N__16195),
            .I(N__16187));
    CascadeMux I__3340 (
            .O(N__16194),
            .I(N__16184));
    CascadeMux I__3339 (
            .O(N__16193),
            .I(N__16181));
    Span4Mux_v I__3338 (
            .O(N__16190),
            .I(N__16176));
    LocalMux I__3337 (
            .O(N__16187),
            .I(N__16176));
    InMux I__3336 (
            .O(N__16184),
            .I(N__16171));
    InMux I__3335 (
            .O(N__16181),
            .I(N__16171));
    Odrv4 I__3334 (
            .O(N__16176),
            .I(measured_delay_hc_17));
    LocalMux I__3333 (
            .O(N__16171),
            .I(measured_delay_hc_17));
    InMux I__3332 (
            .O(N__16166),
            .I(N__16162));
    InMux I__3331 (
            .O(N__16165),
            .I(N__16157));
    LocalMux I__3330 (
            .O(N__16162),
            .I(N__16154));
    InMux I__3329 (
            .O(N__16161),
            .I(N__16149));
    InMux I__3328 (
            .O(N__16160),
            .I(N__16149));
    LocalMux I__3327 (
            .O(N__16157),
            .I(N__16146));
    Span4Mux_v I__3326 (
            .O(N__16154),
            .I(N__16141));
    LocalMux I__3325 (
            .O(N__16149),
            .I(N__16141));
    Odrv12 I__3324 (
            .O(N__16146),
            .I(measured_delay_hc_18));
    Odrv4 I__3323 (
            .O(N__16141),
            .I(measured_delay_hc_18));
    CascadeMux I__3322 (
            .O(N__16136),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_ ));
    InMux I__3321 (
            .O(N__16133),
            .I(N__16127));
    InMux I__3320 (
            .O(N__16132),
            .I(N__16127));
    LocalMux I__3319 (
            .O(N__16127),
            .I(N__16124));
    Span4Mux_h I__3318 (
            .O(N__16124),
            .I(N__16119));
    InMux I__3317 (
            .O(N__16123),
            .I(N__16114));
    InMux I__3316 (
            .O(N__16122),
            .I(N__16114));
    Odrv4 I__3315 (
            .O(N__16119),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    LocalMux I__3314 (
            .O(N__16114),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    CascadeMux I__3313 (
            .O(N__16109),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt8_cascade_ ));
    CascadeMux I__3312 (
            .O(N__16106),
            .I(N__16103));
    InMux I__3311 (
            .O(N__16103),
            .I(N__16098));
    CascadeMux I__3310 (
            .O(N__16102),
            .I(N__16094));
    InMux I__3309 (
            .O(N__16101),
            .I(N__16091));
    LocalMux I__3308 (
            .O(N__16098),
            .I(N__16088));
    CascadeMux I__3307 (
            .O(N__16097),
            .I(N__16085));
    InMux I__3306 (
            .O(N__16094),
            .I(N__16081));
    LocalMux I__3305 (
            .O(N__16091),
            .I(N__16076));
    Span4Mux_v I__3304 (
            .O(N__16088),
            .I(N__16076));
    InMux I__3303 (
            .O(N__16085),
            .I(N__16071));
    InMux I__3302 (
            .O(N__16084),
            .I(N__16071));
    LocalMux I__3301 (
            .O(N__16081),
            .I(measured_delay_hc_8));
    Odrv4 I__3300 (
            .O(N__16076),
            .I(measured_delay_hc_8));
    LocalMux I__3299 (
            .O(N__16071),
            .I(measured_delay_hc_8));
    CascadeMux I__3298 (
            .O(N__16064),
            .I(N__16059));
    InMux I__3297 (
            .O(N__16063),
            .I(N__16056));
    InMux I__3296 (
            .O(N__16062),
            .I(N__16053));
    InMux I__3295 (
            .O(N__16059),
            .I(N__16048));
    LocalMux I__3294 (
            .O(N__16056),
            .I(N__16043));
    LocalMux I__3293 (
            .O(N__16053),
            .I(N__16043));
    InMux I__3292 (
            .O(N__16052),
            .I(N__16038));
    InMux I__3291 (
            .O(N__16051),
            .I(N__16038));
    LocalMux I__3290 (
            .O(N__16048),
            .I(measured_delay_hc_7));
    Odrv12 I__3289 (
            .O(N__16043),
            .I(measured_delay_hc_7));
    LocalMux I__3288 (
            .O(N__16038),
            .I(measured_delay_hc_7));
    CascadeMux I__3287 (
            .O(N__16031),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_ ));
    InMux I__3286 (
            .O(N__16028),
            .I(N__16025));
    LocalMux I__3285 (
            .O(N__16025),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto13 ));
    InMux I__3284 (
            .O(N__16022),
            .I(N__16019));
    LocalMux I__3283 (
            .O(N__16019),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_6 ));
    CascadeMux I__3282 (
            .O(N__16016),
            .I(N__16012));
    InMux I__3281 (
            .O(N__16015),
            .I(N__16006));
    InMux I__3280 (
            .O(N__16012),
            .I(N__16006));
    CascadeMux I__3279 (
            .O(N__16011),
            .I(N__16002));
    LocalMux I__3278 (
            .O(N__16006),
            .I(N__15999));
    InMux I__3277 (
            .O(N__16005),
            .I(N__15994));
    InMux I__3276 (
            .O(N__16002),
            .I(N__15994));
    Span4Mux_v I__3275 (
            .O(N__15999),
            .I(N__15991));
    LocalMux I__3274 (
            .O(N__15994),
            .I(N__15988));
    Odrv4 I__3273 (
            .O(N__15991),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8 ));
    Odrv4 I__3272 (
            .O(N__15988),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8 ));
    CascadeMux I__3271 (
            .O(N__15983),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8_cascade_ ));
    InMux I__3270 (
            .O(N__15980),
            .I(N__15977));
    LocalMux I__3269 (
            .O(N__15977),
            .I(N__15974));
    Span4Mux_v I__3268 (
            .O(N__15974),
            .I(N__15969));
    InMux I__3267 (
            .O(N__15973),
            .I(N__15966));
    InMux I__3266 (
            .O(N__15972),
            .I(N__15963));
    Odrv4 I__3265 (
            .O(N__15969),
            .I(measured_delay_hc_1));
    LocalMux I__3264 (
            .O(N__15966),
            .I(measured_delay_hc_1));
    LocalMux I__3263 (
            .O(N__15963),
            .I(measured_delay_hc_1));
    InMux I__3262 (
            .O(N__15956),
            .I(N__15953));
    LocalMux I__3261 (
            .O(N__15953),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_1 ));
    InMux I__3260 (
            .O(N__15950),
            .I(N__15946));
    InMux I__3259 (
            .O(N__15949),
            .I(N__15943));
    LocalMux I__3258 (
            .O(N__15946),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_2 ));
    LocalMux I__3257 (
            .O(N__15943),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_2 ));
    InMux I__3256 (
            .O(N__15938),
            .I(N__15930));
    InMux I__3255 (
            .O(N__15937),
            .I(N__15930));
    InMux I__3254 (
            .O(N__15936),
            .I(N__15927));
    CascadeMux I__3253 (
            .O(N__15935),
            .I(N__15923));
    LocalMux I__3252 (
            .O(N__15930),
            .I(N__15919));
    LocalMux I__3251 (
            .O(N__15927),
            .I(N__15916));
    InMux I__3250 (
            .O(N__15926),
            .I(N__15913));
    InMux I__3249 (
            .O(N__15923),
            .I(N__15908));
    InMux I__3248 (
            .O(N__15922),
            .I(N__15908));
    Odrv4 I__3247 (
            .O(N__15919),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__3246 (
            .O(N__15916),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3245 (
            .O(N__15913),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3244 (
            .O(N__15908),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__3243 (
            .O(N__15899),
            .I(N__15894));
    CascadeMux I__3242 (
            .O(N__15898),
            .I(N__15891));
    CascadeMux I__3241 (
            .O(N__15897),
            .I(N__15879));
    InMux I__3240 (
            .O(N__15894),
            .I(N__15874));
    InMux I__3239 (
            .O(N__15891),
            .I(N__15874));
    InMux I__3238 (
            .O(N__15890),
            .I(N__15871));
    InMux I__3237 (
            .O(N__15889),
            .I(N__15868));
    InMux I__3236 (
            .O(N__15888),
            .I(N__15855));
    InMux I__3235 (
            .O(N__15887),
            .I(N__15855));
    InMux I__3234 (
            .O(N__15886),
            .I(N__15855));
    InMux I__3233 (
            .O(N__15885),
            .I(N__15855));
    InMux I__3232 (
            .O(N__15884),
            .I(N__15855));
    InMux I__3231 (
            .O(N__15883),
            .I(N__15855));
    InMux I__3230 (
            .O(N__15882),
            .I(N__15846));
    InMux I__3229 (
            .O(N__15879),
            .I(N__15843));
    LocalMux I__3228 (
            .O(N__15874),
            .I(N__15840));
    LocalMux I__3227 (
            .O(N__15871),
            .I(N__15835));
    LocalMux I__3226 (
            .O(N__15868),
            .I(N__15835));
    LocalMux I__3225 (
            .O(N__15855),
            .I(N__15824));
    InMux I__3224 (
            .O(N__15854),
            .I(N__15817));
    InMux I__3223 (
            .O(N__15853),
            .I(N__15817));
    InMux I__3222 (
            .O(N__15852),
            .I(N__15817));
    InMux I__3221 (
            .O(N__15851),
            .I(N__15810));
    InMux I__3220 (
            .O(N__15850),
            .I(N__15810));
    InMux I__3219 (
            .O(N__15849),
            .I(N__15810));
    LocalMux I__3218 (
            .O(N__15846),
            .I(N__15807));
    LocalMux I__3217 (
            .O(N__15843),
            .I(N__15800));
    Span4Mux_v I__3216 (
            .O(N__15840),
            .I(N__15800));
    Span4Mux_v I__3215 (
            .O(N__15835),
            .I(N__15800));
    InMux I__3214 (
            .O(N__15834),
            .I(N__15783));
    InMux I__3213 (
            .O(N__15833),
            .I(N__15783));
    InMux I__3212 (
            .O(N__15832),
            .I(N__15783));
    InMux I__3211 (
            .O(N__15831),
            .I(N__15783));
    InMux I__3210 (
            .O(N__15830),
            .I(N__15783));
    InMux I__3209 (
            .O(N__15829),
            .I(N__15783));
    InMux I__3208 (
            .O(N__15828),
            .I(N__15783));
    InMux I__3207 (
            .O(N__15827),
            .I(N__15783));
    Span4Mux_h I__3206 (
            .O(N__15824),
            .I(N__15778));
    LocalMux I__3205 (
            .O(N__15817),
            .I(N__15778));
    LocalMux I__3204 (
            .O(N__15810),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__3203 (
            .O(N__15807),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__3202 (
            .O(N__15800),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__3201 (
            .O(N__15783),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__3200 (
            .O(N__15778),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__3199 (
            .O(N__15767),
            .I(N__15764));
    InMux I__3198 (
            .O(N__15764),
            .I(N__15756));
    InMux I__3197 (
            .O(N__15763),
            .I(N__15756));
    InMux I__3196 (
            .O(N__15762),
            .I(N__15753));
    InMux I__3195 (
            .O(N__15761),
            .I(N__15750));
    LocalMux I__3194 (
            .O(N__15756),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__3193 (
            .O(N__15753),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__3192 (
            .O(N__15750),
            .I(\phase_controller_inst1.tr_time_passed ));
    CascadeMux I__3191 (
            .O(N__15743),
            .I(N__15725));
    CascadeMux I__3190 (
            .O(N__15742),
            .I(N__15722));
    CascadeMux I__3189 (
            .O(N__15741),
            .I(N__15719));
    CascadeMux I__3188 (
            .O(N__15740),
            .I(N__15716));
    CascadeMux I__3187 (
            .O(N__15739),
            .I(N__15709));
    CascadeMux I__3186 (
            .O(N__15738),
            .I(N__15706));
    CascadeMux I__3185 (
            .O(N__15737),
            .I(N__15703));
    CascadeMux I__3184 (
            .O(N__15736),
            .I(N__15700));
    CascadeMux I__3183 (
            .O(N__15735),
            .I(N__15697));
    CascadeMux I__3182 (
            .O(N__15734),
            .I(N__15694));
    CascadeMux I__3181 (
            .O(N__15733),
            .I(N__15691));
    CascadeMux I__3180 (
            .O(N__15732),
            .I(N__15688));
    InMux I__3179 (
            .O(N__15731),
            .I(N__15669));
    InMux I__3178 (
            .O(N__15730),
            .I(N__15669));
    InMux I__3177 (
            .O(N__15729),
            .I(N__15669));
    InMux I__3176 (
            .O(N__15728),
            .I(N__15669));
    InMux I__3175 (
            .O(N__15725),
            .I(N__15669));
    InMux I__3174 (
            .O(N__15722),
            .I(N__15669));
    InMux I__3173 (
            .O(N__15719),
            .I(N__15669));
    InMux I__3172 (
            .O(N__15716),
            .I(N__15669));
    CascadeMux I__3171 (
            .O(N__15715),
            .I(N__15666));
    InMux I__3170 (
            .O(N__15714),
            .I(N__15657));
    InMux I__3169 (
            .O(N__15713),
            .I(N__15657));
    InMux I__3168 (
            .O(N__15712),
            .I(N__15657));
    InMux I__3167 (
            .O(N__15709),
            .I(N__15657));
    InMux I__3166 (
            .O(N__15706),
            .I(N__15648));
    InMux I__3165 (
            .O(N__15703),
            .I(N__15648));
    InMux I__3164 (
            .O(N__15700),
            .I(N__15648));
    InMux I__3163 (
            .O(N__15697),
            .I(N__15648));
    InMux I__3162 (
            .O(N__15694),
            .I(N__15639));
    InMux I__3161 (
            .O(N__15691),
            .I(N__15639));
    InMux I__3160 (
            .O(N__15688),
            .I(N__15639));
    InMux I__3159 (
            .O(N__15687),
            .I(N__15639));
    CascadeMux I__3158 (
            .O(N__15686),
            .I(N__15636));
    LocalMux I__3157 (
            .O(N__15669),
            .I(N__15633));
    InMux I__3156 (
            .O(N__15666),
            .I(N__15630));
    LocalMux I__3155 (
            .O(N__15657),
            .I(N__15627));
    LocalMux I__3154 (
            .O(N__15648),
            .I(N__15621));
    LocalMux I__3153 (
            .O(N__15639),
            .I(N__15621));
    InMux I__3152 (
            .O(N__15636),
            .I(N__15618));
    Span4Mux_h I__3151 (
            .O(N__15633),
            .I(N__15615));
    LocalMux I__3150 (
            .O(N__15630),
            .I(N__15610));
    Span4Mux_v I__3149 (
            .O(N__15627),
            .I(N__15610));
    InMux I__3148 (
            .O(N__15626),
            .I(N__15607));
    Span4Mux_h I__3147 (
            .O(N__15621),
            .I(N__15604));
    LocalMux I__3146 (
            .O(N__15618),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__3145 (
            .O(N__15615),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__3144 (
            .O(N__15610),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__3143 (
            .O(N__15607),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__3142 (
            .O(N__15604),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__3141 (
            .O(N__15593),
            .I(N__15569));
    InMux I__3140 (
            .O(N__15592),
            .I(N__15569));
    InMux I__3139 (
            .O(N__15591),
            .I(N__15569));
    InMux I__3138 (
            .O(N__15590),
            .I(N__15569));
    InMux I__3137 (
            .O(N__15589),
            .I(N__15569));
    InMux I__3136 (
            .O(N__15588),
            .I(N__15569));
    InMux I__3135 (
            .O(N__15587),
            .I(N__15569));
    InMux I__3134 (
            .O(N__15586),
            .I(N__15569));
    LocalMux I__3133 (
            .O(N__15569),
            .I(N__15563));
    InMux I__3132 (
            .O(N__15568),
            .I(N__15547));
    InMux I__3131 (
            .O(N__15567),
            .I(N__15544));
    InMux I__3130 (
            .O(N__15566),
            .I(N__15541));
    Span4Mux_h I__3129 (
            .O(N__15563),
            .I(N__15538));
    InMux I__3128 (
            .O(N__15562),
            .I(N__15529));
    InMux I__3127 (
            .O(N__15561),
            .I(N__15529));
    InMux I__3126 (
            .O(N__15560),
            .I(N__15529));
    InMux I__3125 (
            .O(N__15559),
            .I(N__15529));
    InMux I__3124 (
            .O(N__15558),
            .I(N__15514));
    InMux I__3123 (
            .O(N__15557),
            .I(N__15514));
    InMux I__3122 (
            .O(N__15556),
            .I(N__15514));
    InMux I__3121 (
            .O(N__15555),
            .I(N__15514));
    InMux I__3120 (
            .O(N__15554),
            .I(N__15514));
    InMux I__3119 (
            .O(N__15553),
            .I(N__15514));
    InMux I__3118 (
            .O(N__15552),
            .I(N__15514));
    InMux I__3117 (
            .O(N__15551),
            .I(N__15511));
    InMux I__3116 (
            .O(N__15550),
            .I(N__15508));
    LocalMux I__3115 (
            .O(N__15547),
            .I(N__15505));
    LocalMux I__3114 (
            .O(N__15544),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__3113 (
            .O(N__15541),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__3112 (
            .O(N__15538),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__3111 (
            .O(N__15529),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__3110 (
            .O(N__15514),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__3109 (
            .O(N__15511),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__3108 (
            .O(N__15508),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__3107 (
            .O(N__15505),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__3106 (
            .O(N__15488),
            .I(N__15485));
    LocalMux I__3105 (
            .O(N__15485),
            .I(\phase_controller_inst1.stoper_tr.N_60 ));
    InMux I__3104 (
            .O(N__15482),
            .I(N__15478));
    InMux I__3103 (
            .O(N__15481),
            .I(N__15474));
    LocalMux I__3102 (
            .O(N__15478),
            .I(N__15471));
    InMux I__3101 (
            .O(N__15477),
            .I(N__15468));
    LocalMux I__3100 (
            .O(N__15474),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__3099 (
            .O(N__15471),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__3098 (
            .O(N__15468),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__3097 (
            .O(N__15461),
            .I(N__15457));
    InMux I__3096 (
            .O(N__15460),
            .I(N__15454));
    LocalMux I__3095 (
            .O(N__15457),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__3094 (
            .O(N__15454),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    IoInMux I__3093 (
            .O(N__15449),
            .I(N__15446));
    LocalMux I__3092 (
            .O(N__15446),
            .I(N__15443));
    Span4Mux_s1_v I__3091 (
            .O(N__15443),
            .I(N__15440));
    Span4Mux_v I__3090 (
            .O(N__15440),
            .I(N__15437));
    Odrv4 I__3089 (
            .O(N__15437),
            .I(\delay_measurement_inst.delay_tr_timer.N_181_i ));
    InMux I__3088 (
            .O(N__15434),
            .I(N__15425));
    InMux I__3087 (
            .O(N__15433),
            .I(N__15425));
    InMux I__3086 (
            .O(N__15432),
            .I(N__15425));
    LocalMux I__3085 (
            .O(N__15425),
            .I(\delay_measurement_inst.hc_prevZ0 ));
    InMux I__3084 (
            .O(N__15422),
            .I(N__15416));
    InMux I__3083 (
            .O(N__15421),
            .I(N__15409));
    InMux I__3082 (
            .O(N__15420),
            .I(N__15409));
    InMux I__3081 (
            .O(N__15419),
            .I(N__15409));
    LocalMux I__3080 (
            .O(N__15416),
            .I(\delay_measurement_inst.hc_syncZ0Z_1 ));
    LocalMux I__3079 (
            .O(N__15409),
            .I(\delay_measurement_inst.hc_syncZ0Z_1 ));
    InMux I__3078 (
            .O(N__15404),
            .I(N__15401));
    LocalMux I__3077 (
            .O(N__15401),
            .I(N__15397));
    InMux I__3076 (
            .O(N__15400),
            .I(N__15394));
    Odrv12 I__3075 (
            .O(N__15397),
            .I(\delay_measurement_inst.delay_hc_timer.N_81 ));
    LocalMux I__3074 (
            .O(N__15394),
            .I(\delay_measurement_inst.delay_hc_timer.N_81 ));
    InMux I__3073 (
            .O(N__15389),
            .I(N__15385));
    InMux I__3072 (
            .O(N__15388),
            .I(N__15382));
    LocalMux I__3071 (
            .O(N__15385),
            .I(N__15378));
    LocalMux I__3070 (
            .O(N__15382),
            .I(N__15375));
    InMux I__3069 (
            .O(N__15381),
            .I(N__15372));
    Odrv4 I__3068 (
            .O(N__15378),
            .I(\delay_measurement_inst.N_54 ));
    Odrv4 I__3067 (
            .O(N__15375),
            .I(\delay_measurement_inst.N_54 ));
    LocalMux I__3066 (
            .O(N__15372),
            .I(\delay_measurement_inst.N_54 ));
    InMux I__3065 (
            .O(N__15365),
            .I(N__15356));
    InMux I__3064 (
            .O(N__15364),
            .I(N__15356));
    InMux I__3063 (
            .O(N__15363),
            .I(N__15349));
    InMux I__3062 (
            .O(N__15362),
            .I(N__15349));
    InMux I__3061 (
            .O(N__15361),
            .I(N__15349));
    LocalMux I__3060 (
            .O(N__15356),
            .I(\delay_measurement_inst.N_132 ));
    LocalMux I__3059 (
            .O(N__15349),
            .I(\delay_measurement_inst.N_132 ));
    CascadeMux I__3058 (
            .O(N__15344),
            .I(N__15340));
    InMux I__3057 (
            .O(N__15343),
            .I(N__15335));
    InMux I__3056 (
            .O(N__15340),
            .I(N__15335));
    LocalMux I__3055 (
            .O(N__15335),
            .I(\delay_measurement_inst.N_139 ));
    CascadeMux I__3054 (
            .O(N__15332),
            .I(N__15329));
    InMux I__3053 (
            .O(N__15329),
            .I(N__15326));
    LocalMux I__3052 (
            .O(N__15326),
            .I(N__15322));
    InMux I__3051 (
            .O(N__15325),
            .I(N__15318));
    Sp12to4 I__3050 (
            .O(N__15322),
            .I(N__15315));
    InMux I__3049 (
            .O(N__15321),
            .I(N__15312));
    LocalMux I__3048 (
            .O(N__15318),
            .I(\delay_measurement_inst.N_134_i ));
    Odrv12 I__3047 (
            .O(N__15315),
            .I(\delay_measurement_inst.N_134_i ));
    LocalMux I__3046 (
            .O(N__15312),
            .I(\delay_measurement_inst.N_134_i ));
    CascadeMux I__3045 (
            .O(N__15305),
            .I(\delay_measurement_inst.N_201_cascade_ ));
    CascadeMux I__3044 (
            .O(N__15302),
            .I(N__15297));
    InMux I__3043 (
            .O(N__15301),
            .I(N__15294));
    InMux I__3042 (
            .O(N__15300),
            .I(N__15289));
    InMux I__3041 (
            .O(N__15297),
            .I(N__15289));
    LocalMux I__3040 (
            .O(N__15294),
            .I(\delay_measurement_inst.delay_tr_timer.N_167 ));
    LocalMux I__3039 (
            .O(N__15289),
            .I(\delay_measurement_inst.delay_tr_timer.N_167 ));
    CascadeMux I__3038 (
            .O(N__15284),
            .I(N__15276));
    CascadeMux I__3037 (
            .O(N__15283),
            .I(N__15273));
    CascadeMux I__3036 (
            .O(N__15282),
            .I(N__15269));
    InMux I__3035 (
            .O(N__15281),
            .I(N__15264));
    InMux I__3034 (
            .O(N__15280),
            .I(N__15264));
    InMux I__3033 (
            .O(N__15279),
            .I(N__15259));
    InMux I__3032 (
            .O(N__15276),
            .I(N__15259));
    InMux I__3031 (
            .O(N__15273),
            .I(N__15252));
    InMux I__3030 (
            .O(N__15272),
            .I(N__15252));
    InMux I__3029 (
            .O(N__15269),
            .I(N__15252));
    LocalMux I__3028 (
            .O(N__15264),
            .I(\delay_measurement_inst.N_170 ));
    LocalMux I__3027 (
            .O(N__15259),
            .I(\delay_measurement_inst.N_170 ));
    LocalMux I__3026 (
            .O(N__15252),
            .I(\delay_measurement_inst.N_170 ));
    CascadeMux I__3025 (
            .O(N__15245),
            .I(N__15240));
    InMux I__3024 (
            .O(N__15244),
            .I(N__15237));
    InMux I__3023 (
            .O(N__15243),
            .I(N__15234));
    InMux I__3022 (
            .O(N__15240),
            .I(N__15231));
    LocalMux I__3021 (
            .O(N__15237),
            .I(N__15226));
    LocalMux I__3020 (
            .O(N__15234),
            .I(N__15226));
    LocalMux I__3019 (
            .O(N__15231),
            .I(N__15223));
    Span4Mux_v I__3018 (
            .O(N__15226),
            .I(N__15220));
    Odrv12 I__3017 (
            .O(N__15223),
            .I(il_min_comp1_D2));
    Odrv4 I__3016 (
            .O(N__15220),
            .I(il_min_comp1_D2));
    InMux I__3015 (
            .O(N__15215),
            .I(N__15211));
    InMux I__3014 (
            .O(N__15214),
            .I(N__15207));
    LocalMux I__3013 (
            .O(N__15211),
            .I(N__15204));
    InMux I__3012 (
            .O(N__15210),
            .I(N__15201));
    LocalMux I__3011 (
            .O(N__15207),
            .I(N__15196));
    Span12Mux_s10_h I__3010 (
            .O(N__15204),
            .I(N__15196));
    LocalMux I__3009 (
            .O(N__15201),
            .I(\phase_controller_inst1.T01_0_sqmuxa ));
    Odrv12 I__3008 (
            .O(N__15196),
            .I(\phase_controller_inst1.T01_0_sqmuxa ));
    InMux I__3007 (
            .O(N__15191),
            .I(N__15186));
    InMux I__3006 (
            .O(N__15190),
            .I(N__15181));
    InMux I__3005 (
            .O(N__15189),
            .I(N__15181));
    LocalMux I__3004 (
            .O(N__15186),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__3003 (
            .O(N__15181),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    IoInMux I__3002 (
            .O(N__15176),
            .I(N__15173));
    LocalMux I__3001 (
            .O(N__15173),
            .I(N__15170));
    Span4Mux_s2_v I__3000 (
            .O(N__15170),
            .I(N__15167));
    Span4Mux_h I__2999 (
            .O(N__15167),
            .I(N__15163));
    CascadeMux I__2998 (
            .O(N__15166),
            .I(N__15160));
    Span4Mux_h I__2997 (
            .O(N__15163),
            .I(N__15157));
    InMux I__2996 (
            .O(N__15160),
            .I(N__15154));
    Odrv4 I__2995 (
            .O(N__15157),
            .I(T12_c));
    LocalMux I__2994 (
            .O(N__15154),
            .I(T12_c));
    InMux I__2993 (
            .O(N__15149),
            .I(N__15146));
    LocalMux I__2992 (
            .O(N__15146),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ));
    CEMux I__2991 (
            .O(N__15143),
            .I(N__15138));
    CEMux I__2990 (
            .O(N__15142),
            .I(N__15135));
    CEMux I__2989 (
            .O(N__15141),
            .I(N__15132));
    LocalMux I__2988 (
            .O(N__15138),
            .I(N__15129));
    LocalMux I__2987 (
            .O(N__15135),
            .I(N__15126));
    LocalMux I__2986 (
            .O(N__15132),
            .I(N__15123));
    Span4Mux_v I__2985 (
            .O(N__15129),
            .I(N__15116));
    Span4Mux_v I__2984 (
            .O(N__15126),
            .I(N__15116));
    Span4Mux_v I__2983 (
            .O(N__15123),
            .I(N__15116));
    Odrv4 I__2982 (
            .O(N__15116),
            .I(\phase_controller_slave.stoper_hc.stoper_state_RNI10KLZ0Z_1 ));
    InMux I__2981 (
            .O(N__15113),
            .I(N__15108));
    CascadeMux I__2980 (
            .O(N__15112),
            .I(N__15104));
    InMux I__2979 (
            .O(N__15111),
            .I(N__15101));
    LocalMux I__2978 (
            .O(N__15108),
            .I(N__15098));
    InMux I__2977 (
            .O(N__15107),
            .I(N__15095));
    InMux I__2976 (
            .O(N__15104),
            .I(N__15092));
    LocalMux I__2975 (
            .O(N__15101),
            .I(N__15089));
    Span4Mux_v I__2974 (
            .O(N__15098),
            .I(N__15082));
    LocalMux I__2973 (
            .O(N__15095),
            .I(N__15082));
    LocalMux I__2972 (
            .O(N__15092),
            .I(N__15082));
    Span4Mux_h I__2971 (
            .O(N__15089),
            .I(N__15079));
    Span4Mux_h I__2970 (
            .O(N__15082),
            .I(N__15076));
    Odrv4 I__2969 (
            .O(N__15079),
            .I(measured_delay_tr_3));
    Odrv4 I__2968 (
            .O(N__15076),
            .I(measured_delay_tr_3));
    InMux I__2967 (
            .O(N__15071),
            .I(N__15068));
    LocalMux I__2966 (
            .O(N__15068),
            .I(N__15063));
    InMux I__2965 (
            .O(N__15067),
            .I(N__15060));
    InMux I__2964 (
            .O(N__15066),
            .I(N__15057));
    Span4Mux_v I__2963 (
            .O(N__15063),
            .I(N__15051));
    LocalMux I__2962 (
            .O(N__15060),
            .I(N__15051));
    LocalMux I__2961 (
            .O(N__15057),
            .I(N__15048));
    InMux I__2960 (
            .O(N__15056),
            .I(N__15045));
    Span4Mux_h I__2959 (
            .O(N__15051),
            .I(N__15042));
    Span12Mux_s5_h I__2958 (
            .O(N__15048),
            .I(N__15037));
    LocalMux I__2957 (
            .O(N__15045),
            .I(N__15037));
    Odrv4 I__2956 (
            .O(N__15042),
            .I(measured_delay_tr_18));
    Odrv12 I__2955 (
            .O(N__15037),
            .I(measured_delay_tr_18));
    InMux I__2954 (
            .O(N__15032),
            .I(N__15029));
    LocalMux I__2953 (
            .O(N__15029),
            .I(N__15025));
    InMux I__2952 (
            .O(N__15028),
            .I(N__15022));
    Span4Mux_v I__2951 (
            .O(N__15025),
            .I(N__15017));
    LocalMux I__2950 (
            .O(N__15022),
            .I(N__15014));
    InMux I__2949 (
            .O(N__15021),
            .I(N__15009));
    InMux I__2948 (
            .O(N__15020),
            .I(N__15009));
    Span4Mux_h I__2947 (
            .O(N__15017),
            .I(N__15004));
    Span4Mux_v I__2946 (
            .O(N__15014),
            .I(N__15004));
    LocalMux I__2945 (
            .O(N__15009),
            .I(N__15001));
    Odrv4 I__2944 (
            .O(N__15004),
            .I(measured_delay_tr_4));
    Odrv4 I__2943 (
            .O(N__15001),
            .I(measured_delay_tr_4));
    InMux I__2942 (
            .O(N__14996),
            .I(N__14992));
    CascadeMux I__2941 (
            .O(N__14995),
            .I(N__14984));
    LocalMux I__2940 (
            .O(N__14992),
            .I(N__14980));
    InMux I__2939 (
            .O(N__14991),
            .I(N__14977));
    InMux I__2938 (
            .O(N__14990),
            .I(N__14970));
    InMux I__2937 (
            .O(N__14989),
            .I(N__14970));
    InMux I__2936 (
            .O(N__14988),
            .I(N__14970));
    InMux I__2935 (
            .O(N__14987),
            .I(N__14963));
    InMux I__2934 (
            .O(N__14984),
            .I(N__14963));
    InMux I__2933 (
            .O(N__14983),
            .I(N__14963));
    Span4Mux_v I__2932 (
            .O(N__14980),
            .I(N__14960));
    LocalMux I__2931 (
            .O(N__14977),
            .I(\delay_measurement_inst.N_129 ));
    LocalMux I__2930 (
            .O(N__14970),
            .I(\delay_measurement_inst.N_129 ));
    LocalMux I__2929 (
            .O(N__14963),
            .I(\delay_measurement_inst.N_129 ));
    Odrv4 I__2928 (
            .O(N__14960),
            .I(\delay_measurement_inst.N_129 ));
    InMux I__2927 (
            .O(N__14951),
            .I(N__14942));
    InMux I__2926 (
            .O(N__14950),
            .I(N__14935));
    InMux I__2925 (
            .O(N__14949),
            .I(N__14935));
    InMux I__2924 (
            .O(N__14948),
            .I(N__14935));
    InMux I__2923 (
            .O(N__14947),
            .I(N__14928));
    InMux I__2922 (
            .O(N__14946),
            .I(N__14928));
    InMux I__2921 (
            .O(N__14945),
            .I(N__14928));
    LocalMux I__2920 (
            .O(N__14942),
            .I(N__14925));
    LocalMux I__2919 (
            .O(N__14935),
            .I(\delay_measurement_inst.N_172 ));
    LocalMux I__2918 (
            .O(N__14928),
            .I(\delay_measurement_inst.N_172 ));
    Odrv4 I__2917 (
            .O(N__14925),
            .I(\delay_measurement_inst.N_172 ));
    InMux I__2916 (
            .O(N__14918),
            .I(N__14915));
    LocalMux I__2915 (
            .O(N__14915),
            .I(N__14911));
    InMux I__2914 (
            .O(N__14914),
            .I(N__14908));
    Span4Mux_h I__2913 (
            .O(N__14911),
            .I(N__14903));
    LocalMux I__2912 (
            .O(N__14908),
            .I(N__14900));
    InMux I__2911 (
            .O(N__14907),
            .I(N__14895));
    InMux I__2910 (
            .O(N__14906),
            .I(N__14895));
    Span4Mux_h I__2909 (
            .O(N__14903),
            .I(N__14892));
    Span4Mux_v I__2908 (
            .O(N__14900),
            .I(N__14887));
    LocalMux I__2907 (
            .O(N__14895),
            .I(N__14887));
    Odrv4 I__2906 (
            .O(N__14892),
            .I(measured_delay_tr_2));
    Odrv4 I__2905 (
            .O(N__14887),
            .I(measured_delay_tr_2));
    CascadeMux I__2904 (
            .O(N__14882),
            .I(N__14878));
    InMux I__2903 (
            .O(N__14881),
            .I(N__14875));
    InMux I__2902 (
            .O(N__14878),
            .I(N__14872));
    LocalMux I__2901 (
            .O(N__14875),
            .I(N__14869));
    LocalMux I__2900 (
            .O(N__14872),
            .I(N__14866));
    Span4Mux_h I__2899 (
            .O(N__14869),
            .I(N__14863));
    Span4Mux_h I__2898 (
            .O(N__14866),
            .I(N__14857));
    Span4Mux_v I__2897 (
            .O(N__14863),
            .I(N__14857));
    InMux I__2896 (
            .O(N__14862),
            .I(N__14854));
    Odrv4 I__2895 (
            .O(N__14857),
            .I(measured_delay_tr_10));
    LocalMux I__2894 (
            .O(N__14854),
            .I(measured_delay_tr_10));
    CascadeMux I__2893 (
            .O(N__14849),
            .I(N__14846));
    InMux I__2892 (
            .O(N__14846),
            .I(N__14843));
    LocalMux I__2891 (
            .O(N__14843),
            .I(N__14838));
    InMux I__2890 (
            .O(N__14842),
            .I(N__14834));
    InMux I__2889 (
            .O(N__14841),
            .I(N__14831));
    Span4Mux_h I__2888 (
            .O(N__14838),
            .I(N__14828));
    InMux I__2887 (
            .O(N__14837),
            .I(N__14825));
    LocalMux I__2886 (
            .O(N__14834),
            .I(N__14822));
    LocalMux I__2885 (
            .O(N__14831),
            .I(N__14819));
    Span4Mux_v I__2884 (
            .O(N__14828),
            .I(N__14814));
    LocalMux I__2883 (
            .O(N__14825),
            .I(N__14814));
    Odrv12 I__2882 (
            .O(N__14822),
            .I(measured_delay_tr_11));
    Odrv4 I__2881 (
            .O(N__14819),
            .I(measured_delay_tr_11));
    Odrv4 I__2880 (
            .O(N__14814),
            .I(measured_delay_tr_11));
    CascadeMux I__2879 (
            .O(N__14807),
            .I(N__14803));
    InMux I__2878 (
            .O(N__14806),
            .I(N__14800));
    InMux I__2877 (
            .O(N__14803),
            .I(N__14797));
    LocalMux I__2876 (
            .O(N__14800),
            .I(N__14794));
    LocalMux I__2875 (
            .O(N__14797),
            .I(N__14791));
    Span4Mux_h I__2874 (
            .O(N__14794),
            .I(N__14788));
    Span4Mux_h I__2873 (
            .O(N__14791),
            .I(N__14784));
    Span4Mux_h I__2872 (
            .O(N__14788),
            .I(N__14781));
    InMux I__2871 (
            .O(N__14787),
            .I(N__14778));
    Odrv4 I__2870 (
            .O(N__14784),
            .I(measured_delay_tr_13));
    Odrv4 I__2869 (
            .O(N__14781),
            .I(measured_delay_tr_13));
    LocalMux I__2868 (
            .O(N__14778),
            .I(measured_delay_tr_13));
    InMux I__2867 (
            .O(N__14771),
            .I(N__14768));
    LocalMux I__2866 (
            .O(N__14768),
            .I(\delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_6 ));
    InMux I__2865 (
            .O(N__14765),
            .I(N__14762));
    LocalMux I__2864 (
            .O(N__14762),
            .I(N__14759));
    Odrv4 I__2863 (
            .O(N__14759),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ));
    InMux I__2862 (
            .O(N__14756),
            .I(N__14753));
    LocalMux I__2861 (
            .O(N__14753),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ));
    InMux I__2860 (
            .O(N__14750),
            .I(N__14747));
    LocalMux I__2859 (
            .O(N__14747),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ));
    InMux I__2858 (
            .O(N__14744),
            .I(N__14741));
    LocalMux I__2857 (
            .O(N__14741),
            .I(N__14738));
    Odrv4 I__2856 (
            .O(N__14738),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ));
    InMux I__2855 (
            .O(N__14735),
            .I(N__14732));
    LocalMux I__2854 (
            .O(N__14732),
            .I(N__14729));
    Odrv4 I__2853 (
            .O(N__14729),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ));
    InMux I__2852 (
            .O(N__14726),
            .I(N__14723));
    LocalMux I__2851 (
            .O(N__14723),
            .I(N__14720));
    Odrv4 I__2850 (
            .O(N__14720),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ));
    InMux I__2849 (
            .O(N__14717),
            .I(N__14714));
    LocalMux I__2848 (
            .O(N__14714),
            .I(N__14711));
    Odrv4 I__2847 (
            .O(N__14711),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ));
    InMux I__2846 (
            .O(N__14708),
            .I(N__14705));
    LocalMux I__2845 (
            .O(N__14705),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ));
    InMux I__2844 (
            .O(N__14702),
            .I(N__14699));
    LocalMux I__2843 (
            .O(N__14699),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__2842 (
            .O(N__14696),
            .I(N__14693));
    InMux I__2841 (
            .O(N__14693),
            .I(N__14690));
    LocalMux I__2840 (
            .O(N__14690),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__2839 (
            .O(N__14687),
            .I(N__14684));
    LocalMux I__2838 (
            .O(N__14684),
            .I(N__14681));
    Span4Mux_h I__2837 (
            .O(N__14681),
            .I(N__14678));
    Odrv4 I__2836 (
            .O(N__14678),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__2835 (
            .O(N__14675),
            .I(N__14672));
    InMux I__2834 (
            .O(N__14672),
            .I(N__14669));
    LocalMux I__2833 (
            .O(N__14669),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    InMux I__2832 (
            .O(N__14666),
            .I(N__14663));
    LocalMux I__2831 (
            .O(N__14663),
            .I(N__14660));
    Odrv4 I__2830 (
            .O(N__14660),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__2829 (
            .O(N__14657),
            .I(N__14654));
    InMux I__2828 (
            .O(N__14654),
            .I(N__14651));
    LocalMux I__2827 (
            .O(N__14651),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    InMux I__2826 (
            .O(N__14648),
            .I(N__14645));
    LocalMux I__2825 (
            .O(N__14645),
            .I(N__14642));
    Odrv4 I__2824 (
            .O(N__14642),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__2823 (
            .O(N__14639),
            .I(N__14636));
    InMux I__2822 (
            .O(N__14636),
            .I(N__14633));
    LocalMux I__2821 (
            .O(N__14633),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    InMux I__2820 (
            .O(N__14630),
            .I(N__14627));
    LocalMux I__2819 (
            .O(N__14627),
            .I(N__14624));
    Odrv4 I__2818 (
            .O(N__14624),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__2817 (
            .O(N__14621),
            .I(N__14618));
    InMux I__2816 (
            .O(N__14618),
            .I(N__14615));
    LocalMux I__2815 (
            .O(N__14615),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__2814 (
            .O(N__14612),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__2813 (
            .O(N__14609),
            .I(N__14606));
    LocalMux I__2812 (
            .O(N__14606),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ));
    InMux I__2811 (
            .O(N__14603),
            .I(N__14600));
    LocalMux I__2810 (
            .O(N__14600),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__2809 (
            .O(N__14597),
            .I(N__14594));
    InMux I__2808 (
            .O(N__14594),
            .I(N__14591));
    LocalMux I__2807 (
            .O(N__14591),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__2806 (
            .O(N__14588),
            .I(N__14585));
    LocalMux I__2805 (
            .O(N__14585),
            .I(N__14582));
    Odrv4 I__2804 (
            .O(N__14582),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__2803 (
            .O(N__14579),
            .I(N__14576));
    InMux I__2802 (
            .O(N__14576),
            .I(N__14573));
    LocalMux I__2801 (
            .O(N__14573),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__2800 (
            .O(N__14570),
            .I(N__14567));
    LocalMux I__2799 (
            .O(N__14567),
            .I(N__14564));
    Odrv4 I__2798 (
            .O(N__14564),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__2797 (
            .O(N__14561),
            .I(N__14558));
    InMux I__2796 (
            .O(N__14558),
            .I(N__14555));
    LocalMux I__2795 (
            .O(N__14555),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__2794 (
            .O(N__14552),
            .I(N__14549));
    InMux I__2793 (
            .O(N__14549),
            .I(N__14546));
    LocalMux I__2792 (
            .O(N__14546),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__2791 (
            .O(N__14543),
            .I(N__14540));
    InMux I__2790 (
            .O(N__14540),
            .I(N__14537));
    LocalMux I__2789 (
            .O(N__14537),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__2788 (
            .O(N__14534),
            .I(N__14531));
    InMux I__2787 (
            .O(N__14531),
            .I(N__14528));
    LocalMux I__2786 (
            .O(N__14528),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__2785 (
            .O(N__14525),
            .I(N__14522));
    InMux I__2784 (
            .O(N__14522),
            .I(N__14519));
    LocalMux I__2783 (
            .O(N__14519),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__2782 (
            .O(N__14516),
            .I(N__14513));
    InMux I__2781 (
            .O(N__14513),
            .I(N__14510));
    LocalMux I__2780 (
            .O(N__14510),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__2779 (
            .O(N__14507),
            .I(N__14504));
    InMux I__2778 (
            .O(N__14504),
            .I(N__14501));
    LocalMux I__2777 (
            .O(N__14501),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__2776 (
            .O(N__14498),
            .I(N__14495));
    LocalMux I__2775 (
            .O(N__14495),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__2774 (
            .O(N__14492),
            .I(N__14489));
    InMux I__2773 (
            .O(N__14489),
            .I(N__14486));
    LocalMux I__2772 (
            .O(N__14486),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__2771 (
            .O(N__14483),
            .I(N__14480));
    LocalMux I__2770 (
            .O(N__14480),
            .I(N__14477));
    Odrv4 I__2769 (
            .O(N__14477),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__2768 (
            .O(N__14474),
            .I(N__14471));
    InMux I__2767 (
            .O(N__14471),
            .I(N__14468));
    LocalMux I__2766 (
            .O(N__14468),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__2765 (
            .O(N__14465),
            .I(N__14462));
    LocalMux I__2764 (
            .O(N__14462),
            .I(N__14459));
    Odrv4 I__2763 (
            .O(N__14459),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__2762 (
            .O(N__14456),
            .I(N__14453));
    InMux I__2761 (
            .O(N__14453),
            .I(N__14450));
    LocalMux I__2760 (
            .O(N__14450),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__2759 (
            .O(N__14447),
            .I(N__14444));
    LocalMux I__2758 (
            .O(N__14444),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__2757 (
            .O(N__14441),
            .I(N__14438));
    InMux I__2756 (
            .O(N__14438),
            .I(N__14435));
    LocalMux I__2755 (
            .O(N__14435),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__2754 (
            .O(N__14432),
            .I(N__14429));
    LocalMux I__2753 (
            .O(N__14429),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__2752 (
            .O(N__14426),
            .I(N__14423));
    InMux I__2751 (
            .O(N__14423),
            .I(N__14420));
    LocalMux I__2750 (
            .O(N__14420),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__2749 (
            .O(N__14417),
            .I(N__14414));
    InMux I__2748 (
            .O(N__14414),
            .I(N__14411));
    LocalMux I__2747 (
            .O(N__14411),
            .I(N__14407));
    InMux I__2746 (
            .O(N__14410),
            .I(N__14404));
    Odrv12 I__2745 (
            .O(N__14407),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    LocalMux I__2744 (
            .O(N__14404),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    CascadeMux I__2743 (
            .O(N__14399),
            .I(N__14394));
    InMux I__2742 (
            .O(N__14398),
            .I(N__14391));
    InMux I__2741 (
            .O(N__14397),
            .I(N__14386));
    InMux I__2740 (
            .O(N__14394),
            .I(N__14386));
    LocalMux I__2739 (
            .O(N__14391),
            .I(N__14383));
    LocalMux I__2738 (
            .O(N__14386),
            .I(N__14380));
    Span4Mux_h I__2737 (
            .O(N__14383),
            .I(N__14377));
    Span4Mux_h I__2736 (
            .O(N__14380),
            .I(N__14374));
    Odrv4 I__2735 (
            .O(N__14377),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    Odrv4 I__2734 (
            .O(N__14374),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    InMux I__2733 (
            .O(N__14369),
            .I(N__14366));
    LocalMux I__2732 (
            .O(N__14366),
            .I(N__14361));
    InMux I__2731 (
            .O(N__14365),
            .I(N__14356));
    InMux I__2730 (
            .O(N__14364),
            .I(N__14356));
    Span4Mux_h I__2729 (
            .O(N__14361),
            .I(N__14353));
    LocalMux I__2728 (
            .O(N__14356),
            .I(N__14350));
    Odrv4 I__2727 (
            .O(N__14353),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    Odrv4 I__2726 (
            .O(N__14350),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    InMux I__2725 (
            .O(N__14345),
            .I(N__14342));
    LocalMux I__2724 (
            .O(N__14342),
            .I(N__14338));
    InMux I__2723 (
            .O(N__14341),
            .I(N__14335));
    Odrv4 I__2722 (
            .O(N__14338),
            .I(\delay_measurement_inst.elapsed_time_hc_6 ));
    LocalMux I__2721 (
            .O(N__14335),
            .I(\delay_measurement_inst.elapsed_time_hc_6 ));
    InMux I__2720 (
            .O(N__14330),
            .I(N__14327));
    LocalMux I__2719 (
            .O(N__14327),
            .I(N__14323));
    CascadeMux I__2718 (
            .O(N__14326),
            .I(N__14320));
    Span4Mux_h I__2717 (
            .O(N__14323),
            .I(N__14317));
    InMux I__2716 (
            .O(N__14320),
            .I(N__14314));
    Span4Mux_h I__2715 (
            .O(N__14317),
            .I(N__14311));
    LocalMux I__2714 (
            .O(N__14314),
            .I(N__14308));
    Odrv4 I__2713 (
            .O(N__14311),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    Odrv4 I__2712 (
            .O(N__14308),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    CascadeMux I__2711 (
            .O(N__14303),
            .I(N__14296));
    InMux I__2710 (
            .O(N__14302),
            .I(N__14287));
    InMux I__2709 (
            .O(N__14301),
            .I(N__14287));
    InMux I__2708 (
            .O(N__14300),
            .I(N__14287));
    InMux I__2707 (
            .O(N__14299),
            .I(N__14287));
    InMux I__2706 (
            .O(N__14296),
            .I(N__14284));
    LocalMux I__2705 (
            .O(N__14287),
            .I(N__14280));
    LocalMux I__2704 (
            .O(N__14284),
            .I(N__14276));
    InMux I__2703 (
            .O(N__14283),
            .I(N__14273));
    Span4Mux_h I__2702 (
            .O(N__14280),
            .I(N__14270));
    InMux I__2701 (
            .O(N__14279),
            .I(N__14267));
    Odrv4 I__2700 (
            .O(N__14276),
            .I(\delay_measurement_inst.N_109 ));
    LocalMux I__2699 (
            .O(N__14273),
            .I(\delay_measurement_inst.N_109 ));
    Odrv4 I__2698 (
            .O(N__14270),
            .I(\delay_measurement_inst.N_109 ));
    LocalMux I__2697 (
            .O(N__14267),
            .I(\delay_measurement_inst.N_109 ));
    InMux I__2696 (
            .O(N__14258),
            .I(N__14242));
    InMux I__2695 (
            .O(N__14257),
            .I(N__14242));
    InMux I__2694 (
            .O(N__14256),
            .I(N__14242));
    InMux I__2693 (
            .O(N__14255),
            .I(N__14242));
    InMux I__2692 (
            .O(N__14254),
            .I(N__14237));
    InMux I__2691 (
            .O(N__14253),
            .I(N__14237));
    InMux I__2690 (
            .O(N__14252),
            .I(N__14232));
    InMux I__2689 (
            .O(N__14251),
            .I(N__14232));
    LocalMux I__2688 (
            .O(N__14242),
            .I(\delay_measurement_inst.N_45 ));
    LocalMux I__2687 (
            .O(N__14237),
            .I(\delay_measurement_inst.N_45 ));
    LocalMux I__2686 (
            .O(N__14232),
            .I(\delay_measurement_inst.N_45 ));
    CascadeMux I__2685 (
            .O(N__14225),
            .I(N__14219));
    CascadeMux I__2684 (
            .O(N__14224),
            .I(N__14216));
    CascadeMux I__2683 (
            .O(N__14223),
            .I(N__14212));
    InMux I__2682 (
            .O(N__14222),
            .I(N__14201));
    InMux I__2681 (
            .O(N__14219),
            .I(N__14201));
    InMux I__2680 (
            .O(N__14216),
            .I(N__14201));
    InMux I__2679 (
            .O(N__14215),
            .I(N__14201));
    InMux I__2678 (
            .O(N__14212),
            .I(N__14196));
    InMux I__2677 (
            .O(N__14211),
            .I(N__14196));
    InMux I__2676 (
            .O(N__14210),
            .I(N__14193));
    LocalMux I__2675 (
            .O(N__14201),
            .I(\delay_measurement_inst.N_107 ));
    LocalMux I__2674 (
            .O(N__14196),
            .I(\delay_measurement_inst.N_107 ));
    LocalMux I__2673 (
            .O(N__14193),
            .I(\delay_measurement_inst.N_107 ));
    InMux I__2672 (
            .O(N__14186),
            .I(N__14183));
    LocalMux I__2671 (
            .O(N__14183),
            .I(N__14179));
    InMux I__2670 (
            .O(N__14182),
            .I(N__14176));
    Odrv4 I__2669 (
            .O(N__14179),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    LocalMux I__2668 (
            .O(N__14176),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    CascadeMux I__2667 (
            .O(N__14171),
            .I(N__14168));
    InMux I__2666 (
            .O(N__14168),
            .I(N__14163));
    InMux I__2665 (
            .O(N__14167),
            .I(N__14158));
    InMux I__2664 (
            .O(N__14166),
            .I(N__14158));
    LocalMux I__2663 (
            .O(N__14163),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__2662 (
            .O(N__14158),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    InMux I__2661 (
            .O(N__14153),
            .I(N__14148));
    InMux I__2660 (
            .O(N__14152),
            .I(N__14143));
    InMux I__2659 (
            .O(N__14151),
            .I(N__14143));
    LocalMux I__2658 (
            .O(N__14148),
            .I(\delay_measurement_inst.tr_prevZ0 ));
    LocalMux I__2657 (
            .O(N__14143),
            .I(\delay_measurement_inst.tr_prevZ0 ));
    CascadeMux I__2656 (
            .O(N__14138),
            .I(N__14134));
    CascadeMux I__2655 (
            .O(N__14137),
            .I(N__14131));
    InMux I__2654 (
            .O(N__14134),
            .I(N__14123));
    InMux I__2653 (
            .O(N__14131),
            .I(N__14123));
    InMux I__2652 (
            .O(N__14130),
            .I(N__14123));
    LocalMux I__2651 (
            .O(N__14123),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    InMux I__2650 (
            .O(N__14120),
            .I(N__14117));
    LocalMux I__2649 (
            .O(N__14117),
            .I(N__14111));
    InMux I__2648 (
            .O(N__14116),
            .I(N__14108));
    InMux I__2647 (
            .O(N__14115),
            .I(N__14103));
    InMux I__2646 (
            .O(N__14114),
            .I(N__14103));
    Span4Mux_h I__2645 (
            .O(N__14111),
            .I(N__14100));
    LocalMux I__2644 (
            .O(N__14108),
            .I(N__14095));
    LocalMux I__2643 (
            .O(N__14103),
            .I(N__14095));
    Odrv4 I__2642 (
            .O(N__14100),
            .I(\delay_measurement_inst.elapsed_time_hc_14 ));
    Odrv4 I__2641 (
            .O(N__14095),
            .I(\delay_measurement_inst.elapsed_time_hc_14 ));
    InMux I__2640 (
            .O(N__14090),
            .I(N__14087));
    LocalMux I__2639 (
            .O(N__14087),
            .I(N__14083));
    CascadeMux I__2638 (
            .O(N__14086),
            .I(N__14079));
    Span4Mux_h I__2637 (
            .O(N__14083),
            .I(N__14076));
    InMux I__2636 (
            .O(N__14082),
            .I(N__14073));
    InMux I__2635 (
            .O(N__14079),
            .I(N__14070));
    Odrv4 I__2634 (
            .O(N__14076),
            .I(\delay_measurement_inst.elapsed_time_hc_9 ));
    LocalMux I__2633 (
            .O(N__14073),
            .I(\delay_measurement_inst.elapsed_time_hc_9 ));
    LocalMux I__2632 (
            .O(N__14070),
            .I(\delay_measurement_inst.elapsed_time_hc_9 ));
    InMux I__2631 (
            .O(N__14063),
            .I(N__14060));
    LocalMux I__2630 (
            .O(N__14060),
            .I(N__14057));
    Span4Mux_h I__2629 (
            .O(N__14057),
            .I(N__14053));
    InMux I__2628 (
            .O(N__14056),
            .I(N__14050));
    Odrv4 I__2627 (
            .O(N__14053),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__2626 (
            .O(N__14050),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    IoInMux I__2625 (
            .O(N__14045),
            .I(N__14042));
    LocalMux I__2624 (
            .O(N__14042),
            .I(N__14038));
    InMux I__2623 (
            .O(N__14041),
            .I(N__14035));
    Span12Mux_s11_v I__2622 (
            .O(N__14038),
            .I(N__14032));
    LocalMux I__2621 (
            .O(N__14035),
            .I(\delay_measurement_inst.delay_hc_timer.N_32 ));
    Odrv12 I__2620 (
            .O(N__14032),
            .I(\delay_measurement_inst.delay_hc_timer.N_32 ));
    InMux I__2619 (
            .O(N__14027),
            .I(N__14018));
    InMux I__2618 (
            .O(N__14026),
            .I(N__14018));
    InMux I__2617 (
            .O(N__14025),
            .I(N__14018));
    LocalMux I__2616 (
            .O(N__14018),
            .I(N__14015));
    Odrv4 I__2615 (
            .O(N__14015),
            .I(\delay_measurement_inst.N_54_i ));
    InMux I__2614 (
            .O(N__14012),
            .I(N__14009));
    LocalMux I__2613 (
            .O(N__14009),
            .I(N__14006));
    Span4Mux_h I__2612 (
            .O(N__14006),
            .I(N__14002));
    InMux I__2611 (
            .O(N__14005),
            .I(N__13999));
    Odrv4 I__2610 (
            .O(N__14002),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__2609 (
            .O(N__13999),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    CascadeMux I__2608 (
            .O(N__13994),
            .I(N__13991));
    InMux I__2607 (
            .O(N__13991),
            .I(N__13988));
    LocalMux I__2606 (
            .O(N__13988),
            .I(N__13985));
    Span4Mux_h I__2605 (
            .O(N__13985),
            .I(N__13982));
    Span4Mux_h I__2604 (
            .O(N__13982),
            .I(N__13979));
    Odrv4 I__2603 (
            .O(N__13979),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    InMux I__2602 (
            .O(N__13976),
            .I(N__13973));
    LocalMux I__2601 (
            .O(N__13973),
            .I(N__13969));
    InMux I__2600 (
            .O(N__13972),
            .I(N__13966));
    Odrv4 I__2599 (
            .O(N__13969),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    LocalMux I__2598 (
            .O(N__13966),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__2597 (
            .O(N__13961),
            .I(N__13958));
    LocalMux I__2596 (
            .O(N__13958),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__2595 (
            .O(N__13955),
            .I(N__13952));
    LocalMux I__2594 (
            .O(N__13952),
            .I(N__13948));
    InMux I__2593 (
            .O(N__13951),
            .I(N__13945));
    Span4Mux_h I__2592 (
            .O(N__13948),
            .I(N__13942));
    LocalMux I__2591 (
            .O(N__13945),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__2590 (
            .O(N__13942),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__2589 (
            .O(N__13937),
            .I(N__13934));
    LocalMux I__2588 (
            .O(N__13934),
            .I(N__13931));
    Span4Mux_s3_v I__2587 (
            .O(N__13931),
            .I(N__13927));
    CascadeMux I__2586 (
            .O(N__13930),
            .I(N__13924));
    Span4Mux_v I__2585 (
            .O(N__13927),
            .I(N__13920));
    InMux I__2584 (
            .O(N__13924),
            .I(N__13917));
    InMux I__2583 (
            .O(N__13923),
            .I(N__13913));
    Span4Mux_v I__2582 (
            .O(N__13920),
            .I(N__13910));
    LocalMux I__2581 (
            .O(N__13917),
            .I(N__13907));
    InMux I__2580 (
            .O(N__13916),
            .I(N__13904));
    LocalMux I__2579 (
            .O(N__13913),
            .I(N__13901));
    Odrv4 I__2578 (
            .O(N__13910),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    Odrv4 I__2577 (
            .O(N__13907),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__2576 (
            .O(N__13904),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    Odrv12 I__2575 (
            .O(N__13901),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    IoInMux I__2574 (
            .O(N__13892),
            .I(N__13889));
    LocalMux I__2573 (
            .O(N__13889),
            .I(s3_phy_c));
    CascadeMux I__2572 (
            .O(N__13886),
            .I(\delay_measurement_inst.N_54_cascade_ ));
    InMux I__2571 (
            .O(N__13883),
            .I(N__13877));
    InMux I__2570 (
            .O(N__13882),
            .I(N__13874));
    InMux I__2569 (
            .O(N__13881),
            .I(N__13869));
    InMux I__2568 (
            .O(N__13880),
            .I(N__13869));
    LocalMux I__2567 (
            .O(N__13877),
            .I(\delay_measurement_inst.tr_syncZ0Z_1 ));
    LocalMux I__2566 (
            .O(N__13874),
            .I(\delay_measurement_inst.tr_syncZ0Z_1 ));
    LocalMux I__2565 (
            .O(N__13869),
            .I(\delay_measurement_inst.tr_syncZ0Z_1 ));
    CascadeMux I__2564 (
            .O(N__13862),
            .I(\delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_5_cascade_ ));
    CascadeMux I__2563 (
            .O(N__13859),
            .I(\delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_9_cascade_ ));
    CascadeMux I__2562 (
            .O(N__13856),
            .I(\delay_measurement_inst.delay_tr_timer.N_160_cascade_ ));
    InMux I__2561 (
            .O(N__13853),
            .I(N__13845));
    InMux I__2560 (
            .O(N__13852),
            .I(N__13845));
    InMux I__2559 (
            .O(N__13851),
            .I(N__13842));
    InMux I__2558 (
            .O(N__13850),
            .I(N__13839));
    LocalMux I__2557 (
            .O(N__13845),
            .I(N__13834));
    LocalMux I__2556 (
            .O(N__13842),
            .I(N__13834));
    LocalMux I__2555 (
            .O(N__13839),
            .I(N__13831));
    Span12Mux_v I__2554 (
            .O(N__13834),
            .I(N__13828));
    Odrv4 I__2553 (
            .O(N__13831),
            .I(\delay_measurement_inst.tr_state_RNIVV8GZ0Z_0 ));
    Odrv12 I__2552 (
            .O(N__13828),
            .I(\delay_measurement_inst.tr_state_RNIVV8GZ0Z_0 ));
    InMux I__2551 (
            .O(N__13823),
            .I(N__13820));
    LocalMux I__2550 (
            .O(N__13820),
            .I(\delay_measurement_inst.delay_tr_timer.un1_reset_i_0 ));
    InMux I__2549 (
            .O(N__13817),
            .I(N__13813));
    InMux I__2548 (
            .O(N__13816),
            .I(N__13810));
    LocalMux I__2547 (
            .O(N__13813),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_2 ));
    LocalMux I__2546 (
            .O(N__13810),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_2 ));
    CascadeMux I__2545 (
            .O(N__13805),
            .I(N__13802));
    InMux I__2544 (
            .O(N__13802),
            .I(N__13799));
    LocalMux I__2543 (
            .O(N__13799),
            .I(N__13795));
    CascadeMux I__2542 (
            .O(N__13798),
            .I(N__13789));
    Span4Mux_h I__2541 (
            .O(N__13795),
            .I(N__13786));
    InMux I__2540 (
            .O(N__13794),
            .I(N__13783));
    InMux I__2539 (
            .O(N__13793),
            .I(N__13780));
    InMux I__2538 (
            .O(N__13792),
            .I(N__13777));
    InMux I__2537 (
            .O(N__13789),
            .I(N__13774));
    Span4Mux_h I__2536 (
            .O(N__13786),
            .I(N__13769));
    LocalMux I__2535 (
            .O(N__13783),
            .I(N__13769));
    LocalMux I__2534 (
            .O(N__13780),
            .I(measured_delay_tr_7));
    LocalMux I__2533 (
            .O(N__13777),
            .I(measured_delay_tr_7));
    LocalMux I__2532 (
            .O(N__13774),
            .I(measured_delay_tr_7));
    Odrv4 I__2531 (
            .O(N__13769),
            .I(measured_delay_tr_7));
    InMux I__2530 (
            .O(N__13760),
            .I(N__13757));
    LocalMux I__2529 (
            .O(N__13757),
            .I(N__13754));
    Span4Mux_h I__2528 (
            .O(N__13754),
            .I(N__13749));
    InMux I__2527 (
            .O(N__13753),
            .I(N__13743));
    InMux I__2526 (
            .O(N__13752),
            .I(N__13743));
    Span4Mux_h I__2525 (
            .O(N__13749),
            .I(N__13740));
    InMux I__2524 (
            .O(N__13748),
            .I(N__13737));
    LocalMux I__2523 (
            .O(N__13743),
            .I(N__13734));
    Odrv4 I__2522 (
            .O(N__13740),
            .I(measured_delay_tr_16));
    LocalMux I__2521 (
            .O(N__13737),
            .I(measured_delay_tr_16));
    Odrv4 I__2520 (
            .O(N__13734),
            .I(measured_delay_tr_16));
    InMux I__2519 (
            .O(N__13727),
            .I(N__13722));
    CascadeMux I__2518 (
            .O(N__13726),
            .I(N__13719));
    InMux I__2517 (
            .O(N__13725),
            .I(N__13715));
    LocalMux I__2516 (
            .O(N__13722),
            .I(N__13709));
    InMux I__2515 (
            .O(N__13719),
            .I(N__13704));
    InMux I__2514 (
            .O(N__13718),
            .I(N__13704));
    LocalMux I__2513 (
            .O(N__13715),
            .I(N__13701));
    InMux I__2512 (
            .O(N__13714),
            .I(N__13698));
    InMux I__2511 (
            .O(N__13713),
            .I(N__13695));
    InMux I__2510 (
            .O(N__13712),
            .I(N__13692));
    Span4Mux_v I__2509 (
            .O(N__13709),
            .I(N__13688));
    LocalMux I__2508 (
            .O(N__13704),
            .I(N__13684));
    Span4Mux_h I__2507 (
            .O(N__13701),
            .I(N__13677));
    LocalMux I__2506 (
            .O(N__13698),
            .I(N__13677));
    LocalMux I__2505 (
            .O(N__13695),
            .I(N__13677));
    LocalMux I__2504 (
            .O(N__13692),
            .I(N__13674));
    InMux I__2503 (
            .O(N__13691),
            .I(N__13671));
    Span4Mux_h I__2502 (
            .O(N__13688),
            .I(N__13668));
    InMux I__2501 (
            .O(N__13687),
            .I(N__13665));
    Span4Mux_h I__2500 (
            .O(N__13684),
            .I(N__13656));
    Span4Mux_v I__2499 (
            .O(N__13677),
            .I(N__13656));
    Span4Mux_v I__2498 (
            .O(N__13674),
            .I(N__13656));
    LocalMux I__2497 (
            .O(N__13671),
            .I(N__13656));
    Odrv4 I__2496 (
            .O(N__13668),
            .I(measured_delay_tr_15));
    LocalMux I__2495 (
            .O(N__13665),
            .I(measured_delay_tr_15));
    Odrv4 I__2494 (
            .O(N__13656),
            .I(measured_delay_tr_15));
    InMux I__2493 (
            .O(N__13649),
            .I(N__13645));
    InMux I__2492 (
            .O(N__13648),
            .I(N__13642));
    LocalMux I__2491 (
            .O(N__13645),
            .I(N__13637));
    LocalMux I__2490 (
            .O(N__13642),
            .I(N__13634));
    InMux I__2489 (
            .O(N__13641),
            .I(N__13629));
    InMux I__2488 (
            .O(N__13640),
            .I(N__13629));
    Span12Mux_v I__2487 (
            .O(N__13637),
            .I(N__13626));
    Span4Mux_h I__2486 (
            .O(N__13634),
            .I(N__13623));
    LocalMux I__2485 (
            .O(N__13629),
            .I(N__13620));
    Odrv12 I__2484 (
            .O(N__13626),
            .I(measured_delay_tr_6));
    Odrv4 I__2483 (
            .O(N__13623),
            .I(measured_delay_tr_6));
    Odrv4 I__2482 (
            .O(N__13620),
            .I(measured_delay_tr_6));
    InMux I__2481 (
            .O(N__13613),
            .I(N__13608));
    InMux I__2480 (
            .O(N__13612),
            .I(N__13605));
    InMux I__2479 (
            .O(N__13611),
            .I(N__13602));
    LocalMux I__2478 (
            .O(N__13608),
            .I(N__13598));
    LocalMux I__2477 (
            .O(N__13605),
            .I(N__13593));
    LocalMux I__2476 (
            .O(N__13602),
            .I(N__13593));
    InMux I__2475 (
            .O(N__13601),
            .I(N__13590));
    Span4Mux_v I__2474 (
            .O(N__13598),
            .I(N__13583));
    Span4Mux_h I__2473 (
            .O(N__13593),
            .I(N__13583));
    LocalMux I__2472 (
            .O(N__13590),
            .I(N__13583));
    Odrv4 I__2471 (
            .O(N__13583),
            .I(measured_delay_tr_12));
    InMux I__2470 (
            .O(N__13580),
            .I(N__13576));
    InMux I__2469 (
            .O(N__13579),
            .I(N__13572));
    LocalMux I__2468 (
            .O(N__13576),
            .I(N__13569));
    InMux I__2467 (
            .O(N__13575),
            .I(N__13566));
    LocalMux I__2466 (
            .O(N__13572),
            .I(N__13563));
    Span4Mux_v I__2465 (
            .O(N__13569),
            .I(N__13558));
    LocalMux I__2464 (
            .O(N__13566),
            .I(N__13558));
    Span4Mux_v I__2463 (
            .O(N__13563),
            .I(N__13552));
    Span4Mux_h I__2462 (
            .O(N__13558),
            .I(N__13552));
    InMux I__2461 (
            .O(N__13557),
            .I(N__13549));
    Odrv4 I__2460 (
            .O(N__13552),
            .I(measured_delay_tr_14));
    LocalMux I__2459 (
            .O(N__13549),
            .I(measured_delay_tr_14));
    CascadeMux I__2458 (
            .O(N__13544),
            .I(N__13541));
    InMux I__2457 (
            .O(N__13541),
            .I(N__13538));
    LocalMux I__2456 (
            .O(N__13538),
            .I(N__13534));
    InMux I__2455 (
            .O(N__13537),
            .I(N__13531));
    Span4Mux_h I__2454 (
            .O(N__13534),
            .I(N__13527));
    LocalMux I__2453 (
            .O(N__13531),
            .I(N__13524));
    InMux I__2452 (
            .O(N__13530),
            .I(N__13521));
    Span4Mux_h I__2451 (
            .O(N__13527),
            .I(N__13518));
    Span4Mux_v I__2450 (
            .O(N__13524),
            .I(N__13513));
    LocalMux I__2449 (
            .O(N__13521),
            .I(N__13513));
    Odrv4 I__2448 (
            .O(N__13518),
            .I(measured_delay_tr_1));
    Odrv4 I__2447 (
            .O(N__13513),
            .I(measured_delay_tr_1));
    InMux I__2446 (
            .O(N__13508),
            .I(N__13505));
    LocalMux I__2445 (
            .O(N__13505),
            .I(N__13500));
    InMux I__2444 (
            .O(N__13504),
            .I(N__13497));
    CascadeMux I__2443 (
            .O(N__13503),
            .I(N__13493));
    Span4Mux_h I__2442 (
            .O(N__13500),
            .I(N__13490));
    LocalMux I__2441 (
            .O(N__13497),
            .I(N__13487));
    InMux I__2440 (
            .O(N__13496),
            .I(N__13484));
    InMux I__2439 (
            .O(N__13493),
            .I(N__13481));
    Odrv4 I__2438 (
            .O(N__13490),
            .I(measured_delay_tr_17));
    Odrv4 I__2437 (
            .O(N__13487),
            .I(measured_delay_tr_17));
    LocalMux I__2436 (
            .O(N__13484),
            .I(measured_delay_tr_17));
    LocalMux I__2435 (
            .O(N__13481),
            .I(measured_delay_tr_17));
    InMux I__2434 (
            .O(N__13472),
            .I(N__13469));
    LocalMux I__2433 (
            .O(N__13469),
            .I(N__13464));
    InMux I__2432 (
            .O(N__13468),
            .I(N__13461));
    InMux I__2431 (
            .O(N__13467),
            .I(N__13458));
    Span4Mux_v I__2430 (
            .O(N__13464),
            .I(N__13453));
    LocalMux I__2429 (
            .O(N__13461),
            .I(N__13450));
    LocalMux I__2428 (
            .O(N__13458),
            .I(N__13447));
    InMux I__2427 (
            .O(N__13457),
            .I(N__13444));
    InMux I__2426 (
            .O(N__13456),
            .I(N__13441));
    Odrv4 I__2425 (
            .O(N__13453),
            .I(measured_delay_tr_9));
    Odrv12 I__2424 (
            .O(N__13450),
            .I(measured_delay_tr_9));
    Odrv4 I__2423 (
            .O(N__13447),
            .I(measured_delay_tr_9));
    LocalMux I__2422 (
            .O(N__13444),
            .I(measured_delay_tr_9));
    LocalMux I__2421 (
            .O(N__13441),
            .I(measured_delay_tr_9));
    InMux I__2420 (
            .O(N__13430),
            .I(N__13427));
    LocalMux I__2419 (
            .O(N__13427),
            .I(N__13423));
    InMux I__2418 (
            .O(N__13426),
            .I(N__13420));
    Span4Mux_v I__2417 (
            .O(N__13423),
            .I(N__13413));
    LocalMux I__2416 (
            .O(N__13420),
            .I(N__13413));
    InMux I__2415 (
            .O(N__13419),
            .I(N__13408));
    InMux I__2414 (
            .O(N__13418),
            .I(N__13408));
    Span4Mux_h I__2413 (
            .O(N__13413),
            .I(N__13405));
    LocalMux I__2412 (
            .O(N__13408),
            .I(N__13402));
    Odrv4 I__2411 (
            .O(N__13405),
            .I(measured_delay_tr_5));
    Odrv4 I__2410 (
            .O(N__13402),
            .I(measured_delay_tr_5));
    InMux I__2409 (
            .O(N__13397),
            .I(N__13393));
    InMux I__2408 (
            .O(N__13396),
            .I(N__13390));
    LocalMux I__2407 (
            .O(N__13393),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__2406 (
            .O(N__13390),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__2405 (
            .O(N__13385),
            .I(N__13382));
    InMux I__2404 (
            .O(N__13382),
            .I(N__13379));
    LocalMux I__2403 (
            .O(N__13379),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ));
    InMux I__2402 (
            .O(N__13376),
            .I(N__13372));
    InMux I__2401 (
            .O(N__13375),
            .I(N__13369));
    LocalMux I__2400 (
            .O(N__13372),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__2399 (
            .O(N__13369),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__2398 (
            .O(N__13364),
            .I(N__13361));
    InMux I__2397 (
            .O(N__13361),
            .I(N__13358));
    LocalMux I__2396 (
            .O(N__13358),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ));
    InMux I__2395 (
            .O(N__13355),
            .I(N__13351));
    InMux I__2394 (
            .O(N__13354),
            .I(N__13348));
    LocalMux I__2393 (
            .O(N__13351),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__2392 (
            .O(N__13348),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__2391 (
            .O(N__13343),
            .I(N__13340));
    InMux I__2390 (
            .O(N__13340),
            .I(N__13337));
    LocalMux I__2389 (
            .O(N__13337),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ));
    InMux I__2388 (
            .O(N__13334),
            .I(N__13330));
    InMux I__2387 (
            .O(N__13333),
            .I(N__13327));
    LocalMux I__2386 (
            .O(N__13330),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__2385 (
            .O(N__13327),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__2384 (
            .O(N__13322),
            .I(N__13319));
    InMux I__2383 (
            .O(N__13319),
            .I(N__13316));
    LocalMux I__2382 (
            .O(N__13316),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ));
    InMux I__2381 (
            .O(N__13313),
            .I(N__13309));
    InMux I__2380 (
            .O(N__13312),
            .I(N__13306));
    LocalMux I__2379 (
            .O(N__13309),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__2378 (
            .O(N__13306),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__2377 (
            .O(N__13301),
            .I(N__13298));
    InMux I__2376 (
            .O(N__13298),
            .I(N__13295));
    LocalMux I__2375 (
            .O(N__13295),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ));
    InMux I__2374 (
            .O(N__13292),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__2373 (
            .O(N__13289),
            .I(N__13278));
    InMux I__2372 (
            .O(N__13288),
            .I(N__13275));
    InMux I__2371 (
            .O(N__13287),
            .I(N__13256));
    InMux I__2370 (
            .O(N__13286),
            .I(N__13256));
    InMux I__2369 (
            .O(N__13285),
            .I(N__13256));
    InMux I__2368 (
            .O(N__13284),
            .I(N__13256));
    InMux I__2367 (
            .O(N__13283),
            .I(N__13256));
    InMux I__2366 (
            .O(N__13282),
            .I(N__13256));
    InMux I__2365 (
            .O(N__13281),
            .I(N__13256));
    InMux I__2364 (
            .O(N__13278),
            .I(N__13245));
    LocalMux I__2363 (
            .O(N__13275),
            .I(N__13242));
    CascadeMux I__2362 (
            .O(N__13274),
            .I(N__13239));
    InMux I__2361 (
            .O(N__13273),
            .I(N__13236));
    CascadeMux I__2360 (
            .O(N__13272),
            .I(N__13233));
    CascadeMux I__2359 (
            .O(N__13271),
            .I(N__13230));
    LocalMux I__2358 (
            .O(N__13256),
            .I(N__13222));
    InMux I__2357 (
            .O(N__13255),
            .I(N__13205));
    InMux I__2356 (
            .O(N__13254),
            .I(N__13205));
    InMux I__2355 (
            .O(N__13253),
            .I(N__13205));
    InMux I__2354 (
            .O(N__13252),
            .I(N__13205));
    InMux I__2353 (
            .O(N__13251),
            .I(N__13205));
    InMux I__2352 (
            .O(N__13250),
            .I(N__13205));
    InMux I__2351 (
            .O(N__13249),
            .I(N__13205));
    InMux I__2350 (
            .O(N__13248),
            .I(N__13205));
    LocalMux I__2349 (
            .O(N__13245),
            .I(N__13202));
    Span4Mux_h I__2348 (
            .O(N__13242),
            .I(N__13199));
    InMux I__2347 (
            .O(N__13239),
            .I(N__13196));
    LocalMux I__2346 (
            .O(N__13236),
            .I(N__13193));
    InMux I__2345 (
            .O(N__13233),
            .I(N__13178));
    InMux I__2344 (
            .O(N__13230),
            .I(N__13178));
    InMux I__2343 (
            .O(N__13229),
            .I(N__13178));
    InMux I__2342 (
            .O(N__13228),
            .I(N__13178));
    InMux I__2341 (
            .O(N__13227),
            .I(N__13178));
    InMux I__2340 (
            .O(N__13226),
            .I(N__13178));
    InMux I__2339 (
            .O(N__13225),
            .I(N__13178));
    Odrv4 I__2338 (
            .O(N__13222),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__2337 (
            .O(N__13205),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__2336 (
            .O(N__13202),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__2335 (
            .O(N__13199),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__2334 (
            .O(N__13196),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__2333 (
            .O(N__13193),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__2332 (
            .O(N__13178),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    InMux I__2331 (
            .O(N__13163),
            .I(N__13158));
    InMux I__2330 (
            .O(N__13162),
            .I(N__13155));
    InMux I__2329 (
            .O(N__13161),
            .I(N__13152));
    LocalMux I__2328 (
            .O(N__13158),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__2327 (
            .O(N__13155),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__2326 (
            .O(N__13152),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__2325 (
            .O(N__13145),
            .I(N__13142));
    LocalMux I__2324 (
            .O(N__13142),
            .I(N__13134));
    InMux I__2323 (
            .O(N__13141),
            .I(N__13131));
    InMux I__2322 (
            .O(N__13140),
            .I(N__13122));
    InMux I__2321 (
            .O(N__13139),
            .I(N__13122));
    InMux I__2320 (
            .O(N__13138),
            .I(N__13122));
    InMux I__2319 (
            .O(N__13137),
            .I(N__13122));
    Odrv12 I__2318 (
            .O(N__13134),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__2317 (
            .O(N__13131),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__2316 (
            .O(N__13122),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__2315 (
            .O(N__13115),
            .I(N__13112));
    InMux I__2314 (
            .O(N__13112),
            .I(N__13109));
    LocalMux I__2313 (
            .O(N__13109),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ));
    InMux I__2312 (
            .O(N__13106),
            .I(N__13103));
    LocalMux I__2311 (
            .O(N__13103),
            .I(N__13100));
    Span12Mux_v I__2310 (
            .O(N__13100),
            .I(N__13097));
    Odrv12 I__2309 (
            .O(N__13097),
            .I(il_min_comp1_D1));
    InMux I__2308 (
            .O(N__13094),
            .I(N__13091));
    LocalMux I__2307 (
            .O(N__13091),
            .I(N__13088));
    Odrv4 I__2306 (
            .O(N__13088),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__2305 (
            .O(N__13085),
            .I(N__13082));
    InMux I__2304 (
            .O(N__13082),
            .I(N__13078));
    InMux I__2303 (
            .O(N__13081),
            .I(N__13075));
    LocalMux I__2302 (
            .O(N__13078),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__2301 (
            .O(N__13075),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__2300 (
            .O(N__13070),
            .I(N__13067));
    InMux I__2299 (
            .O(N__13067),
            .I(N__13064));
    LocalMux I__2298 (
            .O(N__13064),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ));
    InMux I__2297 (
            .O(N__13061),
            .I(N__13057));
    InMux I__2296 (
            .O(N__13060),
            .I(N__13054));
    LocalMux I__2295 (
            .O(N__13057),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__2294 (
            .O(N__13054),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__2293 (
            .O(N__13049),
            .I(N__13046));
    InMux I__2292 (
            .O(N__13046),
            .I(N__13043));
    LocalMux I__2291 (
            .O(N__13043),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ));
    InMux I__2290 (
            .O(N__13040),
            .I(N__13036));
    InMux I__2289 (
            .O(N__13039),
            .I(N__13033));
    LocalMux I__2288 (
            .O(N__13036),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__2287 (
            .O(N__13033),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__2286 (
            .O(N__13028),
            .I(N__13025));
    InMux I__2285 (
            .O(N__13025),
            .I(N__13022));
    LocalMux I__2284 (
            .O(N__13022),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ));
    InMux I__2283 (
            .O(N__13019),
            .I(N__13015));
    InMux I__2282 (
            .O(N__13018),
            .I(N__13012));
    LocalMux I__2281 (
            .O(N__13015),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__2280 (
            .O(N__13012),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__2279 (
            .O(N__13007),
            .I(N__13004));
    InMux I__2278 (
            .O(N__13004),
            .I(N__13001));
    LocalMux I__2277 (
            .O(N__13001),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ));
    InMux I__2276 (
            .O(N__12998),
            .I(N__12994));
    InMux I__2275 (
            .O(N__12997),
            .I(N__12991));
    LocalMux I__2274 (
            .O(N__12994),
            .I(N__12986));
    LocalMux I__2273 (
            .O(N__12991),
            .I(N__12986));
    Span4Mux_h I__2272 (
            .O(N__12986),
            .I(N__12983));
    Odrv4 I__2271 (
            .O(N__12983),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__2270 (
            .O(N__12980),
            .I(N__12977));
    InMux I__2269 (
            .O(N__12977),
            .I(N__12974));
    LocalMux I__2268 (
            .O(N__12974),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ));
    InMux I__2267 (
            .O(N__12971),
            .I(N__12967));
    InMux I__2266 (
            .O(N__12970),
            .I(N__12964));
    LocalMux I__2265 (
            .O(N__12967),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__2264 (
            .O(N__12964),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__2263 (
            .O(N__12959),
            .I(N__12956));
    InMux I__2262 (
            .O(N__12956),
            .I(N__12953));
    LocalMux I__2261 (
            .O(N__12953),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ));
    InMux I__2260 (
            .O(N__12950),
            .I(N__12946));
    InMux I__2259 (
            .O(N__12949),
            .I(N__12943));
    LocalMux I__2258 (
            .O(N__12946),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__2257 (
            .O(N__12943),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__2256 (
            .O(N__12938),
            .I(N__12935));
    InMux I__2255 (
            .O(N__12935),
            .I(N__12932));
    LocalMux I__2254 (
            .O(N__12932),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ));
    InMux I__2253 (
            .O(N__12929),
            .I(N__12926));
    LocalMux I__2252 (
            .O(N__12926),
            .I(N__12923));
    Odrv4 I__2251 (
            .O(N__12923),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__2250 (
            .O(N__12920),
            .I(N__12917));
    InMux I__2249 (
            .O(N__12917),
            .I(N__12914));
    LocalMux I__2248 (
            .O(N__12914),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ));
    InMux I__2247 (
            .O(N__12911),
            .I(N__12908));
    LocalMux I__2246 (
            .O(N__12908),
            .I(N__12905));
    Odrv4 I__2245 (
            .O(N__12905),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ));
    InMux I__2244 (
            .O(N__12902),
            .I(N__12898));
    InMux I__2243 (
            .O(N__12901),
            .I(N__12895));
    LocalMux I__2242 (
            .O(N__12898),
            .I(N__12892));
    LocalMux I__2241 (
            .O(N__12895),
            .I(N__12889));
    Odrv4 I__2240 (
            .O(N__12892),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__2239 (
            .O(N__12889),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__2238 (
            .O(N__12884),
            .I(N__12881));
    InMux I__2237 (
            .O(N__12881),
            .I(N__12878));
    LocalMux I__2236 (
            .O(N__12878),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ));
    InMux I__2235 (
            .O(N__12875),
            .I(N__12872));
    LocalMux I__2234 (
            .O(N__12872),
            .I(N__12869));
    Odrv4 I__2233 (
            .O(N__12869),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ));
    InMux I__2232 (
            .O(N__12866),
            .I(N__12863));
    LocalMux I__2231 (
            .O(N__12863),
            .I(N__12859));
    InMux I__2230 (
            .O(N__12862),
            .I(N__12856));
    Odrv4 I__2229 (
            .O(N__12859),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__2228 (
            .O(N__12856),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__2227 (
            .O(N__12851),
            .I(N__12848));
    InMux I__2226 (
            .O(N__12848),
            .I(N__12845));
    LocalMux I__2225 (
            .O(N__12845),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ));
    InMux I__2224 (
            .O(N__12842),
            .I(N__12839));
    LocalMux I__2223 (
            .O(N__12839),
            .I(N__12836));
    Odrv4 I__2222 (
            .O(N__12836),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ));
    InMux I__2221 (
            .O(N__12833),
            .I(N__12829));
    InMux I__2220 (
            .O(N__12832),
            .I(N__12826));
    LocalMux I__2219 (
            .O(N__12829),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__2218 (
            .O(N__12826),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__2217 (
            .O(N__12821),
            .I(N__12818));
    InMux I__2216 (
            .O(N__12818),
            .I(N__12815));
    LocalMux I__2215 (
            .O(N__12815),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ));
    InMux I__2214 (
            .O(N__12812),
            .I(N__12809));
    LocalMux I__2213 (
            .O(N__12809),
            .I(N__12806));
    Odrv4 I__2212 (
            .O(N__12806),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ));
    InMux I__2211 (
            .O(N__12803),
            .I(N__12799));
    InMux I__2210 (
            .O(N__12802),
            .I(N__12796));
    LocalMux I__2209 (
            .O(N__12799),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__2208 (
            .O(N__12796),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__2207 (
            .O(N__12791),
            .I(N__12788));
    InMux I__2206 (
            .O(N__12788),
            .I(N__12785));
    LocalMux I__2205 (
            .O(N__12785),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ));
    InMux I__2204 (
            .O(N__12782),
            .I(N__12779));
    LocalMux I__2203 (
            .O(N__12779),
            .I(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ));
    CascadeMux I__2202 (
            .O(N__12776),
            .I(N__12773));
    InMux I__2201 (
            .O(N__12773),
            .I(N__12769));
    InMux I__2200 (
            .O(N__12772),
            .I(N__12766));
    LocalMux I__2199 (
            .O(N__12769),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__2198 (
            .O(N__12766),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__2197 (
            .O(N__12761),
            .I(N__12758));
    InMux I__2196 (
            .O(N__12758),
            .I(N__12755));
    LocalMux I__2195 (
            .O(N__12755),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ));
    InMux I__2194 (
            .O(N__12752),
            .I(N__12748));
    InMux I__2193 (
            .O(N__12751),
            .I(N__12745));
    LocalMux I__2192 (
            .O(N__12748),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__2191 (
            .O(N__12745),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__2190 (
            .O(N__12740),
            .I(N__12737));
    InMux I__2189 (
            .O(N__12737),
            .I(N__12734));
    LocalMux I__2188 (
            .O(N__12734),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ));
    InMux I__2187 (
            .O(N__12731),
            .I(N__12728));
    LocalMux I__2186 (
            .O(N__12728),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__2185 (
            .O(N__12725),
            .I(N__12722));
    LocalMux I__2184 (
            .O(N__12722),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_7_9 ));
    CascadeMux I__2183 (
            .O(N__12719),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_6_9_cascade_ ));
    InMux I__2182 (
            .O(N__12716),
            .I(N__12713));
    LocalMux I__2181 (
            .O(N__12713),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ));
    InMux I__2180 (
            .O(N__12710),
            .I(N__12707));
    LocalMux I__2179 (
            .O(N__12707),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__2178 (
            .O(N__12704),
            .I(N__12701));
    LocalMux I__2177 (
            .O(N__12701),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_0_9 ));
    CascadeMux I__2176 (
            .O(N__12698),
            .I(N__12693));
    InMux I__2175 (
            .O(N__12697),
            .I(N__12690));
    InMux I__2174 (
            .O(N__12696),
            .I(N__12687));
    InMux I__2173 (
            .O(N__12693),
            .I(N__12684));
    LocalMux I__2172 (
            .O(N__12690),
            .I(N__12679));
    LocalMux I__2171 (
            .O(N__12687),
            .I(N__12679));
    LocalMux I__2170 (
            .O(N__12684),
            .I(N__12676));
    Odrv4 I__2169 (
            .O(N__12679),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    Odrv4 I__2168 (
            .O(N__12676),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    CascadeMux I__2167 (
            .O(N__12671),
            .I(N__12668));
    InMux I__2166 (
            .O(N__12668),
            .I(N__12663));
    InMux I__2165 (
            .O(N__12667),
            .I(N__12660));
    InMux I__2164 (
            .O(N__12666),
            .I(N__12657));
    LocalMux I__2163 (
            .O(N__12663),
            .I(N__12654));
    LocalMux I__2162 (
            .O(N__12660),
            .I(N__12651));
    LocalMux I__2161 (
            .O(N__12657),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    Odrv4 I__2160 (
            .O(N__12654),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    Odrv4 I__2159 (
            .O(N__12651),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    InMux I__2158 (
            .O(N__12644),
            .I(N__12640));
    InMux I__2157 (
            .O(N__12643),
            .I(N__12637));
    LocalMux I__2156 (
            .O(N__12640),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__2155 (
            .O(N__12637),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    InMux I__2154 (
            .O(N__12632),
            .I(N__12627));
    InMux I__2153 (
            .O(N__12631),
            .I(N__12624));
    InMux I__2152 (
            .O(N__12630),
            .I(N__12620));
    LocalMux I__2151 (
            .O(N__12627),
            .I(N__12615));
    LocalMux I__2150 (
            .O(N__12624),
            .I(N__12615));
    InMux I__2149 (
            .O(N__12623),
            .I(N__12612));
    LocalMux I__2148 (
            .O(N__12620),
            .I(N__12608));
    Span4Mux_v I__2147 (
            .O(N__12615),
            .I(N__12603));
    LocalMux I__2146 (
            .O(N__12612),
            .I(N__12603));
    InMux I__2145 (
            .O(N__12611),
            .I(N__12600));
    Span12Mux_v I__2144 (
            .O(N__12608),
            .I(N__12597));
    Span4Mux_v I__2143 (
            .O(N__12603),
            .I(N__12594));
    LocalMux I__2142 (
            .O(N__12600),
            .I(measured_delay_tr_8));
    Odrv12 I__2141 (
            .O(N__12597),
            .I(measured_delay_tr_8));
    Odrv4 I__2140 (
            .O(N__12594),
            .I(measured_delay_tr_8));
    InMux I__2139 (
            .O(N__12587),
            .I(N__12584));
    LocalMux I__2138 (
            .O(N__12584),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__2137 (
            .O(N__12581),
            .I(N__12578));
    LocalMux I__2136 (
            .O(N__12578),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    CascadeMux I__2135 (
            .O(N__12575),
            .I(N__12572));
    InMux I__2134 (
            .O(N__12572),
            .I(N__12569));
    LocalMux I__2133 (
            .O(N__12569),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__2132 (
            .O(N__12566),
            .I(N__12563));
    LocalMux I__2131 (
            .O(N__12563),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__2130 (
            .O(N__12560),
            .I(N__12557));
    LocalMux I__2129 (
            .O(N__12557),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__2128 (
            .O(N__12554),
            .I(N__12551));
    LocalMux I__2127 (
            .O(N__12551),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    CascadeMux I__2126 (
            .O(N__12548),
            .I(N__12545));
    InMux I__2125 (
            .O(N__12545),
            .I(N__12542));
    LocalMux I__2124 (
            .O(N__12542),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__2123 (
            .O(N__12539),
            .I(N__12536));
    LocalMux I__2122 (
            .O(N__12536),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__2121 (
            .O(N__12533),
            .I(N__12530));
    LocalMux I__2120 (
            .O(N__12530),
            .I(\delay_measurement_inst.delay_hc_timer.N_101 ));
    CascadeMux I__2119 (
            .O(N__12527),
            .I(\delay_measurement_inst.delay_hc_timer.N_81_cascade_ ));
    InMux I__2118 (
            .O(N__12524),
            .I(N__12521));
    LocalMux I__2117 (
            .O(N__12521),
            .I(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_4 ));
    CascadeMux I__2116 (
            .O(N__12518),
            .I(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_6_cascade_ ));
    InMux I__2115 (
            .O(N__12515),
            .I(N__12512));
    LocalMux I__2114 (
            .O(N__12512),
            .I(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_5 ));
    InMux I__2113 (
            .O(N__12509),
            .I(N__12503));
    InMux I__2112 (
            .O(N__12508),
            .I(N__12503));
    LocalMux I__2111 (
            .O(N__12503),
            .I(\delay_measurement_inst.delay_hc_timer.N_105 ));
    InMux I__2110 (
            .O(N__12500),
            .I(N__12497));
    LocalMux I__2109 (
            .O(N__12497),
            .I(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_0 ));
    CascadeMux I__2108 (
            .O(N__12494),
            .I(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_9_cascade_ ));
    InMux I__2107 (
            .O(N__12491),
            .I(N__12488));
    LocalMux I__2106 (
            .O(N__12488),
            .I(N__12484));
    InMux I__2105 (
            .O(N__12487),
            .I(N__12481));
    Span4Mux_v I__2104 (
            .O(N__12484),
            .I(N__12476));
    LocalMux I__2103 (
            .O(N__12481),
            .I(N__12476));
    Odrv4 I__2102 (
            .O(N__12476),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    InMux I__2101 (
            .O(N__12473),
            .I(N__12469));
    InMux I__2100 (
            .O(N__12472),
            .I(N__12466));
    LocalMux I__2099 (
            .O(N__12469),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__2098 (
            .O(N__12466),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__2097 (
            .O(N__12461),
            .I(N__12458));
    LocalMux I__2096 (
            .O(N__12458),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__2095 (
            .O(N__12455),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__2094 (
            .O(N__12452),
            .I(N__12448));
    InMux I__2093 (
            .O(N__12451),
            .I(N__12445));
    LocalMux I__2092 (
            .O(N__12448),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__2091 (
            .O(N__12445),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__2090 (
            .O(N__12440),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__2089 (
            .O(N__12437),
            .I(N__12434));
    LocalMux I__2088 (
            .O(N__12434),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    IoInMux I__2087 (
            .O(N__12431),
            .I(N__12428));
    LocalMux I__2086 (
            .O(N__12428),
            .I(N__12425));
    Span4Mux_s3_v I__2085 (
            .O(N__12425),
            .I(N__12422));
    Sp12to4 I__2084 (
            .O(N__12422),
            .I(N__12419));
    Span12Mux_s9_h I__2083 (
            .O(N__12419),
            .I(N__12416));
    Span12Mux_v I__2082 (
            .O(N__12416),
            .I(N__12413));
    Odrv12 I__2081 (
            .O(N__12413),
            .I(\delay_measurement_inst.delay_tr_timer.N_180_i ));
    InMux I__2080 (
            .O(N__12410),
            .I(N__12407));
    LocalMux I__2079 (
            .O(N__12407),
            .I(N__12404));
    Odrv12 I__2078 (
            .O(N__12404),
            .I(il_min_comp1_c));
    InMux I__2077 (
            .O(N__12401),
            .I(N__12398));
    LocalMux I__2076 (
            .O(N__12398),
            .I(N__12394));
    InMux I__2075 (
            .O(N__12397),
            .I(N__12391));
    Odrv4 I__2074 (
            .O(N__12394),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__2073 (
            .O(N__12391),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__2072 (
            .O(N__12386),
            .I(N__12383));
    InMux I__2071 (
            .O(N__12383),
            .I(N__12380));
    LocalMux I__2070 (
            .O(N__12380),
            .I(N__12377));
    Odrv4 I__2069 (
            .O(N__12377),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__2068 (
            .O(N__12374),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__2067 (
            .O(N__12371),
            .I(N__12367));
    InMux I__2066 (
            .O(N__12370),
            .I(N__12364));
    LocalMux I__2065 (
            .O(N__12367),
            .I(N__12361));
    LocalMux I__2064 (
            .O(N__12364),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__2063 (
            .O(N__12361),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__2062 (
            .O(N__12356),
            .I(N__12353));
    LocalMux I__2061 (
            .O(N__12353),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__2060 (
            .O(N__12350),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__2059 (
            .O(N__12347),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__2058 (
            .O(N__12344),
            .I(N__12340));
    InMux I__2057 (
            .O(N__12343),
            .I(N__12337));
    LocalMux I__2056 (
            .O(N__12340),
            .I(N__12334));
    LocalMux I__2055 (
            .O(N__12337),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__2054 (
            .O(N__12334),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__2053 (
            .O(N__12329),
            .I(N__12326));
    LocalMux I__2052 (
            .O(N__12326),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__2051 (
            .O(N__12323),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    CascadeMux I__2050 (
            .O(N__12320),
            .I(N__12316));
    InMux I__2049 (
            .O(N__12319),
            .I(N__12313));
    InMux I__2048 (
            .O(N__12316),
            .I(N__12310));
    LocalMux I__2047 (
            .O(N__12313),
            .I(N__12307));
    LocalMux I__2046 (
            .O(N__12310),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__2045 (
            .O(N__12307),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__2044 (
            .O(N__12302),
            .I(N__12299));
    InMux I__2043 (
            .O(N__12299),
            .I(N__12296));
    LocalMux I__2042 (
            .O(N__12296),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__2041 (
            .O(N__12293),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__2040 (
            .O(N__12290),
            .I(N__12286));
    InMux I__2039 (
            .O(N__12289),
            .I(N__12283));
    LocalMux I__2038 (
            .O(N__12286),
            .I(N__12280));
    LocalMux I__2037 (
            .O(N__12283),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__2036 (
            .O(N__12280),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__2035 (
            .O(N__12275),
            .I(N__12272));
    LocalMux I__2034 (
            .O(N__12272),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    InMux I__2033 (
            .O(N__12269),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__2032 (
            .O(N__12266),
            .I(N__12262));
    InMux I__2031 (
            .O(N__12265),
            .I(N__12259));
    LocalMux I__2030 (
            .O(N__12262),
            .I(N__12256));
    LocalMux I__2029 (
            .O(N__12259),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__2028 (
            .O(N__12256),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__2027 (
            .O(N__12251),
            .I(N__12248));
    InMux I__2026 (
            .O(N__12248),
            .I(N__12245));
    LocalMux I__2025 (
            .O(N__12245),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__2024 (
            .O(N__12242),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__2023 (
            .O(N__12239),
            .I(N__12235));
    InMux I__2022 (
            .O(N__12238),
            .I(N__12232));
    LocalMux I__2021 (
            .O(N__12235),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__2020 (
            .O(N__12232),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__2019 (
            .O(N__12227),
            .I(N__12224));
    LocalMux I__2018 (
            .O(N__12224),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    InMux I__2017 (
            .O(N__12221),
            .I(bfn_8_27_0_));
    InMux I__2016 (
            .O(N__12218),
            .I(N__12215));
    LocalMux I__2015 (
            .O(N__12215),
            .I(N__12212));
    Odrv4 I__2014 (
            .O(N__12212),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    InMux I__2013 (
            .O(N__12209),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__2012 (
            .O(N__12206),
            .I(N__12202));
    InMux I__2011 (
            .O(N__12205),
            .I(N__12199));
    LocalMux I__2010 (
            .O(N__12202),
            .I(N__12196));
    LocalMux I__2009 (
            .O(N__12199),
            .I(N__12193));
    Odrv4 I__2008 (
            .O(N__12196),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__2007 (
            .O(N__12193),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__2006 (
            .O(N__12188),
            .I(N__12185));
    InMux I__2005 (
            .O(N__12185),
            .I(N__12182));
    LocalMux I__2004 (
            .O(N__12182),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0 ));
    InMux I__2003 (
            .O(N__12179),
            .I(N__12176));
    LocalMux I__2002 (
            .O(N__12176),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    InMux I__2001 (
            .O(N__12173),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__2000 (
            .O(N__12170),
            .I(N__12166));
    InMux I__1999 (
            .O(N__12169),
            .I(N__12163));
    LocalMux I__1998 (
            .O(N__12166),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__1997 (
            .O(N__12163),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__1996 (
            .O(N__12158),
            .I(N__12155));
    LocalMux I__1995 (
            .O(N__12155),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__1994 (
            .O(N__12152),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__1993 (
            .O(N__12149),
            .I(N__12145));
    InMux I__1992 (
            .O(N__12148),
            .I(N__12142));
    LocalMux I__1991 (
            .O(N__12145),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__1990 (
            .O(N__12142),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__1989 (
            .O(N__12137),
            .I(N__12134));
    LocalMux I__1988 (
            .O(N__12134),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__1987 (
            .O(N__12131),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__1986 (
            .O(N__12128),
            .I(N__12124));
    InMux I__1985 (
            .O(N__12127),
            .I(N__12121));
    LocalMux I__1984 (
            .O(N__12124),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__1983 (
            .O(N__12121),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__1982 (
            .O(N__12116),
            .I(N__12113));
    LocalMux I__1981 (
            .O(N__12113),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__1980 (
            .O(N__12110),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__1979 (
            .O(N__12107),
            .I(N__12103));
    InMux I__1978 (
            .O(N__12106),
            .I(N__12100));
    LocalMux I__1977 (
            .O(N__12103),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__1976 (
            .O(N__12100),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__1975 (
            .O(N__12095),
            .I(N__12092));
    LocalMux I__1974 (
            .O(N__12092),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__1973 (
            .O(N__12089),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__1972 (
            .O(N__12086),
            .I(N__12083));
    LocalMux I__1971 (
            .O(N__12083),
            .I(N__12079));
    InMux I__1970 (
            .O(N__12082),
            .I(N__12076));
    Odrv4 I__1969 (
            .O(N__12079),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__1968 (
            .O(N__12076),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__1967 (
            .O(N__12071),
            .I(N__12068));
    LocalMux I__1966 (
            .O(N__12068),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    InMux I__1965 (
            .O(N__12065),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__1964 (
            .O(N__12062),
            .I(N__12059));
    LocalMux I__1963 (
            .O(N__12059),
            .I(N__12055));
    InMux I__1962 (
            .O(N__12058),
            .I(N__12052));
    Odrv4 I__1961 (
            .O(N__12055),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__1960 (
            .O(N__12052),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__1959 (
            .O(N__12047),
            .I(N__12044));
    LocalMux I__1958 (
            .O(N__12044),
            .I(N__12041));
    Odrv4 I__1957 (
            .O(N__12041),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    InMux I__1956 (
            .O(N__12038),
            .I(bfn_8_26_0_));
    CEMux I__1955 (
            .O(N__12035),
            .I(N__12032));
    LocalMux I__1954 (
            .O(N__12032),
            .I(N__12026));
    CEMux I__1953 (
            .O(N__12031),
            .I(N__12023));
    CEMux I__1952 (
            .O(N__12030),
            .I(N__12020));
    CEMux I__1951 (
            .O(N__12029),
            .I(N__12017));
    Span4Mux_v I__1950 (
            .O(N__12026),
            .I(N__12011));
    LocalMux I__1949 (
            .O(N__12023),
            .I(N__12011));
    LocalMux I__1948 (
            .O(N__12020),
            .I(N__12008));
    LocalMux I__1947 (
            .O(N__12017),
            .I(N__12005));
    CEMux I__1946 (
            .O(N__12016),
            .I(N__12002));
    Span4Mux_h I__1945 (
            .O(N__12011),
            .I(N__11999));
    Span4Mux_v I__1944 (
            .O(N__12008),
            .I(N__11994));
    Span4Mux_h I__1943 (
            .O(N__12005),
            .I(N__11994));
    LocalMux I__1942 (
            .O(N__12002),
            .I(N__11991));
    Odrv4 I__1941 (
            .O(N__11999),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1 ));
    Odrv4 I__1940 (
            .O(N__11994),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1 ));
    Odrv12 I__1939 (
            .O(N__11991),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1 ));
    CascadeMux I__1938 (
            .O(N__11984),
            .I(N__11981));
    InMux I__1937 (
            .O(N__11981),
            .I(N__11977));
    InMux I__1936 (
            .O(N__11980),
            .I(N__11974));
    LocalMux I__1935 (
            .O(N__11977),
            .I(N__11968));
    LocalMux I__1934 (
            .O(N__11974),
            .I(N__11968));
    InMux I__1933 (
            .O(N__11973),
            .I(N__11965));
    Odrv4 I__1932 (
            .O(N__11968),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__1931 (
            .O(N__11965),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__1930 (
            .O(N__11960),
            .I(N__11957));
    InMux I__1929 (
            .O(N__11957),
            .I(N__11954));
    LocalMux I__1928 (
            .O(N__11954),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    InMux I__1927 (
            .O(N__11951),
            .I(N__11948));
    LocalMux I__1926 (
            .O(N__11948),
            .I(N__11944));
    InMux I__1925 (
            .O(N__11947),
            .I(N__11941));
    Odrv4 I__1924 (
            .O(N__11944),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__1923 (
            .O(N__11941),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__1922 (
            .O(N__11936),
            .I(N__11933));
    LocalMux I__1921 (
            .O(N__11933),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__1920 (
            .O(N__11930),
            .I(N__11927));
    LocalMux I__1919 (
            .O(N__11927),
            .I(N__11924));
    Span4Mux_h I__1918 (
            .O(N__11924),
            .I(N__11921));
    Odrv4 I__1917 (
            .O(N__11921),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__1916 (
            .O(N__11918),
            .I(N__11915));
    LocalMux I__1915 (
            .O(N__11915),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    InMux I__1914 (
            .O(N__11912),
            .I(N__11909));
    LocalMux I__1913 (
            .O(N__11909),
            .I(N__11906));
    Sp12to4 I__1912 (
            .O(N__11906),
            .I(N__11903));
    Odrv12 I__1911 (
            .O(N__11903),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__1910 (
            .O(N__11900),
            .I(N__11894));
    InMux I__1909 (
            .O(N__11899),
            .I(N__11883));
    InMux I__1908 (
            .O(N__11898),
            .I(N__11883));
    InMux I__1907 (
            .O(N__11897),
            .I(N__11883));
    InMux I__1906 (
            .O(N__11894),
            .I(N__11878));
    InMux I__1905 (
            .O(N__11893),
            .I(N__11878));
    CascadeMux I__1904 (
            .O(N__11892),
            .I(N__11869));
    InMux I__1903 (
            .O(N__11891),
            .I(N__11864));
    InMux I__1902 (
            .O(N__11890),
            .I(N__11864));
    LocalMux I__1901 (
            .O(N__11883),
            .I(N__11861));
    LocalMux I__1900 (
            .O(N__11878),
            .I(N__11858));
    InMux I__1899 (
            .O(N__11877),
            .I(N__11847));
    InMux I__1898 (
            .O(N__11876),
            .I(N__11847));
    InMux I__1897 (
            .O(N__11875),
            .I(N__11847));
    InMux I__1896 (
            .O(N__11874),
            .I(N__11847));
    InMux I__1895 (
            .O(N__11873),
            .I(N__11847));
    CascadeMux I__1894 (
            .O(N__11872),
            .I(N__11844));
    InMux I__1893 (
            .O(N__11869),
            .I(N__11835));
    LocalMux I__1892 (
            .O(N__11864),
            .I(N__11832));
    Span4Mux_v I__1891 (
            .O(N__11861),
            .I(N__11825));
    Span4Mux_v I__1890 (
            .O(N__11858),
            .I(N__11825));
    LocalMux I__1889 (
            .O(N__11847),
            .I(N__11825));
    InMux I__1888 (
            .O(N__11844),
            .I(N__11818));
    InMux I__1887 (
            .O(N__11843),
            .I(N__11818));
    InMux I__1886 (
            .O(N__11842),
            .I(N__11818));
    InMux I__1885 (
            .O(N__11841),
            .I(N__11811));
    InMux I__1884 (
            .O(N__11840),
            .I(N__11811));
    InMux I__1883 (
            .O(N__11839),
            .I(N__11811));
    InMux I__1882 (
            .O(N__11838),
            .I(N__11808));
    LocalMux I__1881 (
            .O(N__11835),
            .I(N__11803));
    Span4Mux_h I__1880 (
            .O(N__11832),
            .I(N__11803));
    Span4Mux_h I__1879 (
            .O(N__11825),
            .I(N__11800));
    LocalMux I__1878 (
            .O(N__11818),
            .I(\phase_controller_inst1.stoper_tr.un3_start ));
    LocalMux I__1877 (
            .O(N__11811),
            .I(\phase_controller_inst1.stoper_tr.un3_start ));
    LocalMux I__1876 (
            .O(N__11808),
            .I(\phase_controller_inst1.stoper_tr.un3_start ));
    Odrv4 I__1875 (
            .O(N__11803),
            .I(\phase_controller_inst1.stoper_tr.un3_start ));
    Odrv4 I__1874 (
            .O(N__11800),
            .I(\phase_controller_inst1.stoper_tr.un3_start ));
    CascadeMux I__1873 (
            .O(N__11789),
            .I(N__11778));
    CascadeMux I__1872 (
            .O(N__11788),
            .I(N__11774));
    CascadeMux I__1871 (
            .O(N__11787),
            .I(N__11771));
    CascadeMux I__1870 (
            .O(N__11786),
            .I(N__11767));
    CascadeMux I__1869 (
            .O(N__11785),
            .I(N__11764));
    CascadeMux I__1868 (
            .O(N__11784),
            .I(N__11758));
    CascadeMux I__1867 (
            .O(N__11783),
            .I(N__11755));
    CascadeMux I__1866 (
            .O(N__11782),
            .I(N__11752));
    InMux I__1865 (
            .O(N__11781),
            .I(N__11742));
    InMux I__1864 (
            .O(N__11778),
            .I(N__11735));
    InMux I__1863 (
            .O(N__11777),
            .I(N__11735));
    InMux I__1862 (
            .O(N__11774),
            .I(N__11735));
    InMux I__1861 (
            .O(N__11771),
            .I(N__11724));
    InMux I__1860 (
            .O(N__11770),
            .I(N__11724));
    InMux I__1859 (
            .O(N__11767),
            .I(N__11724));
    InMux I__1858 (
            .O(N__11764),
            .I(N__11724));
    InMux I__1857 (
            .O(N__11763),
            .I(N__11724));
    InMux I__1856 (
            .O(N__11762),
            .I(N__11717));
    InMux I__1855 (
            .O(N__11761),
            .I(N__11717));
    InMux I__1854 (
            .O(N__11758),
            .I(N__11717));
    InMux I__1853 (
            .O(N__11755),
            .I(N__11708));
    InMux I__1852 (
            .O(N__11752),
            .I(N__11708));
    InMux I__1851 (
            .O(N__11751),
            .I(N__11708));
    InMux I__1850 (
            .O(N__11750),
            .I(N__11708));
    CascadeMux I__1849 (
            .O(N__11749),
            .I(N__11703));
    CascadeMux I__1848 (
            .O(N__11748),
            .I(N__11698));
    CascadeMux I__1847 (
            .O(N__11747),
            .I(N__11695));
    CascadeMux I__1846 (
            .O(N__11746),
            .I(N__11692));
    CascadeMux I__1845 (
            .O(N__11745),
            .I(N__11689));
    LocalMux I__1844 (
            .O(N__11742),
            .I(N__11686));
    LocalMux I__1843 (
            .O(N__11735),
            .I(N__11683));
    LocalMux I__1842 (
            .O(N__11724),
            .I(N__11676));
    LocalMux I__1841 (
            .O(N__11717),
            .I(N__11676));
    LocalMux I__1840 (
            .O(N__11708),
            .I(N__11676));
    InMux I__1839 (
            .O(N__11707),
            .I(N__11670));
    InMux I__1838 (
            .O(N__11706),
            .I(N__11667));
    InMux I__1837 (
            .O(N__11703),
            .I(N__11658));
    InMux I__1836 (
            .O(N__11702),
            .I(N__11658));
    InMux I__1835 (
            .O(N__11701),
            .I(N__11658));
    InMux I__1834 (
            .O(N__11698),
            .I(N__11658));
    InMux I__1833 (
            .O(N__11695),
            .I(N__11651));
    InMux I__1832 (
            .O(N__11692),
            .I(N__11651));
    InMux I__1831 (
            .O(N__11689),
            .I(N__11651));
    Span4Mux_v I__1830 (
            .O(N__11686),
            .I(N__11644));
    Span4Mux_v I__1829 (
            .O(N__11683),
            .I(N__11644));
    Span4Mux_v I__1828 (
            .O(N__11676),
            .I(N__11644));
    InMux I__1827 (
            .O(N__11675),
            .I(N__11639));
    InMux I__1826 (
            .O(N__11674),
            .I(N__11639));
    InMux I__1825 (
            .O(N__11673),
            .I(N__11636));
    LocalMux I__1824 (
            .O(N__11670),
            .I(N__11633));
    LocalMux I__1823 (
            .O(N__11667),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2 ));
    LocalMux I__1822 (
            .O(N__11658),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2 ));
    LocalMux I__1821 (
            .O(N__11651),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2 ));
    Odrv4 I__1820 (
            .O(N__11644),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2 ));
    LocalMux I__1819 (
            .O(N__11639),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2 ));
    LocalMux I__1818 (
            .O(N__11636),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2 ));
    Odrv4 I__1817 (
            .O(N__11633),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2 ));
    InMux I__1816 (
            .O(N__11618),
            .I(N__11602));
    InMux I__1815 (
            .O(N__11617),
            .I(N__11602));
    InMux I__1814 (
            .O(N__11616),
            .I(N__11602));
    InMux I__1813 (
            .O(N__11615),
            .I(N__11591));
    InMux I__1812 (
            .O(N__11614),
            .I(N__11591));
    InMux I__1811 (
            .O(N__11613),
            .I(N__11591));
    InMux I__1810 (
            .O(N__11612),
            .I(N__11591));
    InMux I__1809 (
            .O(N__11611),
            .I(N__11591));
    InMux I__1808 (
            .O(N__11610),
            .I(N__11586));
    InMux I__1807 (
            .O(N__11609),
            .I(N__11586));
    LocalMux I__1806 (
            .O(N__11602),
            .I(N__11572));
    LocalMux I__1805 (
            .O(N__11591),
            .I(N__11567));
    LocalMux I__1804 (
            .O(N__11586),
            .I(N__11567));
    InMux I__1803 (
            .O(N__11585),
            .I(N__11560));
    InMux I__1802 (
            .O(N__11584),
            .I(N__11560));
    InMux I__1801 (
            .O(N__11583),
            .I(N__11560));
    InMux I__1800 (
            .O(N__11582),
            .I(N__11551));
    InMux I__1799 (
            .O(N__11581),
            .I(N__11551));
    InMux I__1798 (
            .O(N__11580),
            .I(N__11551));
    InMux I__1797 (
            .O(N__11579),
            .I(N__11551));
    InMux I__1796 (
            .O(N__11578),
            .I(N__11542));
    InMux I__1795 (
            .O(N__11577),
            .I(N__11542));
    InMux I__1794 (
            .O(N__11576),
            .I(N__11542));
    InMux I__1793 (
            .O(N__11575),
            .I(N__11542));
    Span4Mux_v I__1792 (
            .O(N__11572),
            .I(N__11535));
    Span4Mux_v I__1791 (
            .O(N__11567),
            .I(N__11535));
    LocalMux I__1790 (
            .O(N__11560),
            .I(N__11532));
    LocalMux I__1789 (
            .O(N__11551),
            .I(N__11529));
    LocalMux I__1788 (
            .O(N__11542),
            .I(N__11526));
    InMux I__1787 (
            .O(N__11541),
            .I(N__11523));
    InMux I__1786 (
            .O(N__11540),
            .I(N__11520));
    Odrv4 I__1785 (
            .O(N__11535),
            .I(\phase_controller_inst1.stoper_tr.un1_startlt15 ));
    Odrv4 I__1784 (
            .O(N__11532),
            .I(\phase_controller_inst1.stoper_tr.un1_startlt15 ));
    Odrv12 I__1783 (
            .O(N__11529),
            .I(\phase_controller_inst1.stoper_tr.un1_startlt15 ));
    Odrv4 I__1782 (
            .O(N__11526),
            .I(\phase_controller_inst1.stoper_tr.un1_startlt15 ));
    LocalMux I__1781 (
            .O(N__11523),
            .I(\phase_controller_inst1.stoper_tr.un1_startlt15 ));
    LocalMux I__1780 (
            .O(N__11520),
            .I(\phase_controller_inst1.stoper_tr.un1_startlt15 ));
    InMux I__1779 (
            .O(N__11507),
            .I(N__11504));
    LocalMux I__1778 (
            .O(N__11504),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__1777 (
            .O(N__11501),
            .I(N__11498));
    InMux I__1776 (
            .O(N__11498),
            .I(N__11495));
    LocalMux I__1775 (
            .O(N__11495),
            .I(N__11492));
    Odrv4 I__1774 (
            .O(N__11492),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ));
    InMux I__1773 (
            .O(N__11489),
            .I(N__11486));
    LocalMux I__1772 (
            .O(N__11486),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__1771 (
            .O(N__11483),
            .I(N__11480));
    LocalMux I__1770 (
            .O(N__11480),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ));
    InMux I__1769 (
            .O(N__11477),
            .I(N__11441));
    InMux I__1768 (
            .O(N__11476),
            .I(N__11441));
    InMux I__1767 (
            .O(N__11475),
            .I(N__11441));
    InMux I__1766 (
            .O(N__11474),
            .I(N__11441));
    InMux I__1765 (
            .O(N__11473),
            .I(N__11441));
    InMux I__1764 (
            .O(N__11472),
            .I(N__11441));
    InMux I__1763 (
            .O(N__11471),
            .I(N__11441));
    InMux I__1762 (
            .O(N__11470),
            .I(N__11441));
    InMux I__1761 (
            .O(N__11469),
            .I(N__11430));
    InMux I__1760 (
            .O(N__11468),
            .I(N__11430));
    InMux I__1759 (
            .O(N__11467),
            .I(N__11430));
    InMux I__1758 (
            .O(N__11466),
            .I(N__11430));
    InMux I__1757 (
            .O(N__11465),
            .I(N__11430));
    InMux I__1756 (
            .O(N__11464),
            .I(N__11411));
    InMux I__1755 (
            .O(N__11463),
            .I(N__11411));
    InMux I__1754 (
            .O(N__11462),
            .I(N__11411));
    InMux I__1753 (
            .O(N__11461),
            .I(N__11411));
    InMux I__1752 (
            .O(N__11460),
            .I(N__11411));
    InMux I__1751 (
            .O(N__11459),
            .I(N__11411));
    InMux I__1750 (
            .O(N__11458),
            .I(N__11411));
    LocalMux I__1749 (
            .O(N__11441),
            .I(N__11406));
    LocalMux I__1748 (
            .O(N__11430),
            .I(N__11406));
    InMux I__1747 (
            .O(N__11429),
            .I(N__11403));
    InMux I__1746 (
            .O(N__11428),
            .I(N__11400));
    InMux I__1745 (
            .O(N__11427),
            .I(N__11397));
    InMux I__1744 (
            .O(N__11426),
            .I(N__11394));
    LocalMux I__1743 (
            .O(N__11411),
            .I(N__11387));
    Span4Mux_v I__1742 (
            .O(N__11406),
            .I(N__11387));
    LocalMux I__1741 (
            .O(N__11403),
            .I(N__11387));
    LocalMux I__1740 (
            .O(N__11400),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    LocalMux I__1739 (
            .O(N__11397),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    LocalMux I__1738 (
            .O(N__11394),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__1737 (
            .O(N__11387),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    CascadeMux I__1736 (
            .O(N__11378),
            .I(N__11375));
    InMux I__1735 (
            .O(N__11375),
            .I(N__11372));
    LocalMux I__1734 (
            .O(N__11372),
            .I(N__11369));
    Odrv4 I__1733 (
            .O(N__11369),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ));
    CascadeMux I__1732 (
            .O(N__11366),
            .I(N__11353));
    CascadeMux I__1731 (
            .O(N__11365),
            .I(N__11347));
    CascadeMux I__1730 (
            .O(N__11364),
            .I(N__11344));
    CascadeMux I__1729 (
            .O(N__11363),
            .I(N__11341));
    CascadeMux I__1728 (
            .O(N__11362),
            .I(N__11338));
    CascadeMux I__1727 (
            .O(N__11361),
            .I(N__11334));
    InMux I__1726 (
            .O(N__11360),
            .I(N__11326));
    InMux I__1725 (
            .O(N__11359),
            .I(N__11326));
    CascadeMux I__1724 (
            .O(N__11358),
            .I(N__11319));
    CascadeMux I__1723 (
            .O(N__11357),
            .I(N__11316));
    CascadeMux I__1722 (
            .O(N__11356),
            .I(N__11313));
    InMux I__1721 (
            .O(N__11353),
            .I(N__11309));
    InMux I__1720 (
            .O(N__11352),
            .I(N__11294));
    InMux I__1719 (
            .O(N__11351),
            .I(N__11294));
    InMux I__1718 (
            .O(N__11350),
            .I(N__11294));
    InMux I__1717 (
            .O(N__11347),
            .I(N__11294));
    InMux I__1716 (
            .O(N__11344),
            .I(N__11294));
    InMux I__1715 (
            .O(N__11341),
            .I(N__11294));
    InMux I__1714 (
            .O(N__11338),
            .I(N__11294));
    InMux I__1713 (
            .O(N__11337),
            .I(N__11283));
    InMux I__1712 (
            .O(N__11334),
            .I(N__11283));
    InMux I__1711 (
            .O(N__11333),
            .I(N__11283));
    InMux I__1710 (
            .O(N__11332),
            .I(N__11283));
    InMux I__1709 (
            .O(N__11331),
            .I(N__11283));
    LocalMux I__1708 (
            .O(N__11326),
            .I(N__11280));
    InMux I__1707 (
            .O(N__11325),
            .I(N__11263));
    InMux I__1706 (
            .O(N__11324),
            .I(N__11263));
    InMux I__1705 (
            .O(N__11323),
            .I(N__11263));
    InMux I__1704 (
            .O(N__11322),
            .I(N__11263));
    InMux I__1703 (
            .O(N__11319),
            .I(N__11263));
    InMux I__1702 (
            .O(N__11316),
            .I(N__11263));
    InMux I__1701 (
            .O(N__11313),
            .I(N__11263));
    InMux I__1700 (
            .O(N__11312),
            .I(N__11263));
    LocalMux I__1699 (
            .O(N__11309),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1698 (
            .O(N__11294),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1697 (
            .O(N__11283),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__1696 (
            .O(N__11280),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1695 (
            .O(N__11263),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__1694 (
            .O(N__11252),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto9_cZ0_cascade_ ));
    InMux I__1693 (
            .O(N__11249),
            .I(N__11246));
    LocalMux I__1692 (
            .O(N__11246),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto13 ));
    CascadeMux I__1691 (
            .O(N__11243),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_6_cascade_ ));
    CascadeMux I__1690 (
            .O(N__11240),
            .I(N__11236));
    InMux I__1689 (
            .O(N__11239),
            .I(N__11231));
    InMux I__1688 (
            .O(N__11236),
            .I(N__11231));
    LocalMux I__1687 (
            .O(N__11231),
            .I(N__11227));
    CascadeMux I__1686 (
            .O(N__11230),
            .I(N__11223));
    Span4Mux_h I__1685 (
            .O(N__11227),
            .I(N__11220));
    InMux I__1684 (
            .O(N__11226),
            .I(N__11215));
    InMux I__1683 (
            .O(N__11223),
            .I(N__11215));
    Odrv4 I__1682 (
            .O(N__11220),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8 ));
    LocalMux I__1681 (
            .O(N__11215),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8 ));
    CascadeMux I__1680 (
            .O(N__11210),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8_cascade_ ));
    CascadeMux I__1679 (
            .O(N__11207),
            .I(N__11203));
    CascadeMux I__1678 (
            .O(N__11206),
            .I(N__11199));
    InMux I__1677 (
            .O(N__11203),
            .I(N__11195));
    InMux I__1676 (
            .O(N__11202),
            .I(N__11192));
    InMux I__1675 (
            .O(N__11199),
            .I(N__11187));
    InMux I__1674 (
            .O(N__11198),
            .I(N__11187));
    LocalMux I__1673 (
            .O(N__11195),
            .I(N__11182));
    LocalMux I__1672 (
            .O(N__11192),
            .I(N__11182));
    LocalMux I__1671 (
            .O(N__11187),
            .I(N__11176));
    Span4Mux_h I__1670 (
            .O(N__11182),
            .I(N__11176));
    InMux I__1669 (
            .O(N__11181),
            .I(N__11173));
    Odrv4 I__1668 (
            .O(N__11176),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_9 ));
    LocalMux I__1667 (
            .O(N__11173),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_9 ));
    CascadeMux I__1666 (
            .O(N__11168),
            .I(N__11165));
    InMux I__1665 (
            .O(N__11165),
            .I(N__11162));
    LocalMux I__1664 (
            .O(N__11162),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DKZ0 ));
    CascadeMux I__1663 (
            .O(N__11159),
            .I(N__11156));
    InMux I__1662 (
            .O(N__11156),
            .I(N__11153));
    LocalMux I__1661 (
            .O(N__11153),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__1660 (
            .O(N__11150),
            .I(N__11147));
    LocalMux I__1659 (
            .O(N__11147),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ));
    InMux I__1658 (
            .O(N__11144),
            .I(N__11141));
    LocalMux I__1657 (
            .O(N__11141),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ));
    CascadeMux I__1656 (
            .O(N__11138),
            .I(N__11135));
    InMux I__1655 (
            .O(N__11135),
            .I(N__11132));
    LocalMux I__1654 (
            .O(N__11132),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ));
    InMux I__1653 (
            .O(N__11129),
            .I(N__11126));
    LocalMux I__1652 (
            .O(N__11126),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ));
    CascadeMux I__1651 (
            .O(N__11123),
            .I(N__11120));
    InMux I__1650 (
            .O(N__11120),
            .I(N__11117));
    LocalMux I__1649 (
            .O(N__11117),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ));
    InMux I__1648 (
            .O(N__11114),
            .I(N__11111));
    LocalMux I__1647 (
            .O(N__11111),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__1646 (
            .O(N__11108),
            .I(N__11105));
    LocalMux I__1645 (
            .O(N__11105),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ));
    CascadeMux I__1644 (
            .O(N__11102),
            .I(N__11099));
    InMux I__1643 (
            .O(N__11099),
            .I(N__11096));
    LocalMux I__1642 (
            .O(N__11096),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ));
    InMux I__1641 (
            .O(N__11093),
            .I(N__11090));
    LocalMux I__1640 (
            .O(N__11090),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ));
    CascadeMux I__1639 (
            .O(N__11087),
            .I(N__11084));
    InMux I__1638 (
            .O(N__11084),
            .I(N__11081));
    LocalMux I__1637 (
            .O(N__11081),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ));
    InMux I__1636 (
            .O(N__11078),
            .I(N__11075));
    LocalMux I__1635 (
            .O(N__11075),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ));
    CascadeMux I__1634 (
            .O(N__11072),
            .I(N__11069));
    InMux I__1633 (
            .O(N__11069),
            .I(N__11066));
    LocalMux I__1632 (
            .O(N__11066),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ));
    CascadeMux I__1631 (
            .O(N__11063),
            .I(N__11060));
    InMux I__1630 (
            .O(N__11060),
            .I(N__11057));
    LocalMux I__1629 (
            .O(N__11057),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    CascadeMux I__1628 (
            .O(N__11054),
            .I(N__11049));
    CascadeMux I__1627 (
            .O(N__11053),
            .I(N__11046));
    InMux I__1626 (
            .O(N__11052),
            .I(N__11043));
    InMux I__1625 (
            .O(N__11049),
            .I(N__11038));
    InMux I__1624 (
            .O(N__11046),
            .I(N__11038));
    LocalMux I__1623 (
            .O(N__11043),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__1622 (
            .O(N__11038),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__1621 (
            .O(N__11033),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__1620 (
            .O(N__11030),
            .I(N__11025));
    CascadeMux I__1619 (
            .O(N__11029),
            .I(N__11022));
    InMux I__1618 (
            .O(N__11028),
            .I(N__11019));
    InMux I__1617 (
            .O(N__11025),
            .I(N__11014));
    InMux I__1616 (
            .O(N__11022),
            .I(N__11014));
    LocalMux I__1615 (
            .O(N__11019),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__1614 (
            .O(N__11014),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__1613 (
            .O(N__11009),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__1612 (
            .O(N__11006),
            .I(N__11001));
    InMux I__1611 (
            .O(N__11005),
            .I(N__10998));
    InMux I__1610 (
            .O(N__11004),
            .I(N__10995));
    LocalMux I__1609 (
            .O(N__11001),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__1608 (
            .O(N__10998),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__1607 (
            .O(N__10995),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__1606 (
            .O(N__10988),
            .I(bfn_8_16_0_));
    InMux I__1605 (
            .O(N__10985),
            .I(N__10980));
    InMux I__1604 (
            .O(N__10984),
            .I(N__10977));
    InMux I__1603 (
            .O(N__10983),
            .I(N__10974));
    LocalMux I__1602 (
            .O(N__10980),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__1601 (
            .O(N__10977),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__1600 (
            .O(N__10974),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__1599 (
            .O(N__10967),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__1598 (
            .O(N__10964),
            .I(N__10960));
    InMux I__1597 (
            .O(N__10963),
            .I(N__10957));
    LocalMux I__1596 (
            .O(N__10960),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__1595 (
            .O(N__10957),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    CascadeMux I__1594 (
            .O(N__10952),
            .I(N__10947));
    CascadeMux I__1593 (
            .O(N__10951),
            .I(N__10944));
    InMux I__1592 (
            .O(N__10950),
            .I(N__10941));
    InMux I__1591 (
            .O(N__10947),
            .I(N__10936));
    InMux I__1590 (
            .O(N__10944),
            .I(N__10936));
    LocalMux I__1589 (
            .O(N__10941),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__1588 (
            .O(N__10936),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__1587 (
            .O(N__10931),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__1586 (
            .O(N__10928),
            .I(N__10924));
    InMux I__1585 (
            .O(N__10927),
            .I(N__10921));
    LocalMux I__1584 (
            .O(N__10924),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__1583 (
            .O(N__10921),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__1582 (
            .O(N__10916),
            .I(N__10911));
    CascadeMux I__1581 (
            .O(N__10915),
            .I(N__10908));
    InMux I__1580 (
            .O(N__10914),
            .I(N__10905));
    InMux I__1579 (
            .O(N__10911),
            .I(N__10900));
    InMux I__1578 (
            .O(N__10908),
            .I(N__10900));
    LocalMux I__1577 (
            .O(N__10905),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__1576 (
            .O(N__10900),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__1575 (
            .O(N__10895),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__1574 (
            .O(N__10892),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__1573 (
            .O(N__10889),
            .I(N__10874));
    CEMux I__1572 (
            .O(N__10888),
            .I(N__10874));
    CEMux I__1571 (
            .O(N__10887),
            .I(N__10874));
    CEMux I__1570 (
            .O(N__10886),
            .I(N__10874));
    CEMux I__1569 (
            .O(N__10885),
            .I(N__10874));
    GlobalMux I__1568 (
            .O(N__10874),
            .I(N__10871));
    gio2CtrlBuf I__1567 (
            .O(N__10871),
            .I(\delay_measurement_inst.delay_hc_timer.N_178_i_g ));
    CascadeMux I__1566 (
            .O(N__10868),
            .I(N__10865));
    InMux I__1565 (
            .O(N__10865),
            .I(N__10862));
    LocalMux I__1564 (
            .O(N__10862),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ));
    InMux I__1563 (
            .O(N__10859),
            .I(N__10854));
    InMux I__1562 (
            .O(N__10858),
            .I(N__10849));
    InMux I__1561 (
            .O(N__10857),
            .I(N__10849));
    LocalMux I__1560 (
            .O(N__10854),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__1559 (
            .O(N__10849),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__1558 (
            .O(N__10844),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__1557 (
            .O(N__10841),
            .I(N__10836));
    CascadeMux I__1556 (
            .O(N__10840),
            .I(N__10833));
    InMux I__1555 (
            .O(N__10839),
            .I(N__10830));
    InMux I__1554 (
            .O(N__10836),
            .I(N__10825));
    InMux I__1553 (
            .O(N__10833),
            .I(N__10825));
    LocalMux I__1552 (
            .O(N__10830),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__1551 (
            .O(N__10825),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__1550 (
            .O(N__10820),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__1549 (
            .O(N__10817),
            .I(N__10812));
    CascadeMux I__1548 (
            .O(N__10816),
            .I(N__10809));
    InMux I__1547 (
            .O(N__10815),
            .I(N__10806));
    InMux I__1546 (
            .O(N__10812),
            .I(N__10801));
    InMux I__1545 (
            .O(N__10809),
            .I(N__10801));
    LocalMux I__1544 (
            .O(N__10806),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__1543 (
            .O(N__10801),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__1542 (
            .O(N__10796),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__1541 (
            .O(N__10793),
            .I(N__10788));
    InMux I__1540 (
            .O(N__10792),
            .I(N__10785));
    InMux I__1539 (
            .O(N__10791),
            .I(N__10782));
    LocalMux I__1538 (
            .O(N__10788),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__1537 (
            .O(N__10785),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__1536 (
            .O(N__10782),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__1535 (
            .O(N__10775),
            .I(bfn_8_15_0_));
    InMux I__1534 (
            .O(N__10772),
            .I(N__10767));
    InMux I__1533 (
            .O(N__10771),
            .I(N__10764));
    InMux I__1532 (
            .O(N__10770),
            .I(N__10761));
    LocalMux I__1531 (
            .O(N__10767),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__1530 (
            .O(N__10764),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__1529 (
            .O(N__10761),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__1528 (
            .O(N__10754),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__1527 (
            .O(N__10751),
            .I(N__10746));
    CascadeMux I__1526 (
            .O(N__10750),
            .I(N__10743));
    InMux I__1525 (
            .O(N__10749),
            .I(N__10740));
    InMux I__1524 (
            .O(N__10746),
            .I(N__10735));
    InMux I__1523 (
            .O(N__10743),
            .I(N__10735));
    LocalMux I__1522 (
            .O(N__10740),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__1521 (
            .O(N__10735),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__1520 (
            .O(N__10730),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__1519 (
            .O(N__10727),
            .I(N__10722));
    CascadeMux I__1518 (
            .O(N__10726),
            .I(N__10719));
    InMux I__1517 (
            .O(N__10725),
            .I(N__10716));
    InMux I__1516 (
            .O(N__10722),
            .I(N__10711));
    InMux I__1515 (
            .O(N__10719),
            .I(N__10711));
    LocalMux I__1514 (
            .O(N__10716),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__1513 (
            .O(N__10711),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__1512 (
            .O(N__10706),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__1511 (
            .O(N__10703),
            .I(N__10698));
    InMux I__1510 (
            .O(N__10702),
            .I(N__10693));
    InMux I__1509 (
            .O(N__10701),
            .I(N__10693));
    LocalMux I__1508 (
            .O(N__10698),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__1507 (
            .O(N__10693),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__1506 (
            .O(N__10688),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__1505 (
            .O(N__10685),
            .I(N__10680));
    InMux I__1504 (
            .O(N__10684),
            .I(N__10675));
    InMux I__1503 (
            .O(N__10683),
            .I(N__10675));
    LocalMux I__1502 (
            .O(N__10680),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__1501 (
            .O(N__10675),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__1500 (
            .O(N__10670),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__1499 (
            .O(N__10667),
            .I(N__10662));
    InMux I__1498 (
            .O(N__10666),
            .I(N__10657));
    InMux I__1497 (
            .O(N__10665),
            .I(N__10657));
    LocalMux I__1496 (
            .O(N__10662),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__1495 (
            .O(N__10657),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__1494 (
            .O(N__10652),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__1493 (
            .O(N__10649),
            .I(N__10644));
    CascadeMux I__1492 (
            .O(N__10648),
            .I(N__10641));
    InMux I__1491 (
            .O(N__10647),
            .I(N__10638));
    InMux I__1490 (
            .O(N__10644),
            .I(N__10633));
    InMux I__1489 (
            .O(N__10641),
            .I(N__10633));
    LocalMux I__1488 (
            .O(N__10638),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__1487 (
            .O(N__10633),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__1486 (
            .O(N__10628),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__1485 (
            .O(N__10625),
            .I(N__10620));
    CascadeMux I__1484 (
            .O(N__10624),
            .I(N__10617));
    InMux I__1483 (
            .O(N__10623),
            .I(N__10614));
    InMux I__1482 (
            .O(N__10620),
            .I(N__10609));
    InMux I__1481 (
            .O(N__10617),
            .I(N__10609));
    LocalMux I__1480 (
            .O(N__10614),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__1479 (
            .O(N__10609),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__1478 (
            .O(N__10604),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__1477 (
            .O(N__10601),
            .I(N__10596));
    InMux I__1476 (
            .O(N__10600),
            .I(N__10593));
    InMux I__1475 (
            .O(N__10599),
            .I(N__10590));
    LocalMux I__1474 (
            .O(N__10596),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__1473 (
            .O(N__10593),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__1472 (
            .O(N__10590),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__1471 (
            .O(N__10583),
            .I(bfn_8_14_0_));
    InMux I__1470 (
            .O(N__10580),
            .I(N__10575));
    InMux I__1469 (
            .O(N__10579),
            .I(N__10572));
    InMux I__1468 (
            .O(N__10578),
            .I(N__10569));
    LocalMux I__1467 (
            .O(N__10575),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__1466 (
            .O(N__10572),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__1465 (
            .O(N__10569),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__1464 (
            .O(N__10562),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__1463 (
            .O(N__10559),
            .I(N__10554));
    CascadeMux I__1462 (
            .O(N__10558),
            .I(N__10551));
    InMux I__1461 (
            .O(N__10557),
            .I(N__10548));
    InMux I__1460 (
            .O(N__10554),
            .I(N__10543));
    InMux I__1459 (
            .O(N__10551),
            .I(N__10543));
    LocalMux I__1458 (
            .O(N__10548),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__1457 (
            .O(N__10543),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__1456 (
            .O(N__10538),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__1455 (
            .O(N__10535),
            .I(N__10530));
    CascadeMux I__1454 (
            .O(N__10534),
            .I(N__10527));
    InMux I__1453 (
            .O(N__10533),
            .I(N__10524));
    InMux I__1452 (
            .O(N__10530),
            .I(N__10519));
    InMux I__1451 (
            .O(N__10527),
            .I(N__10519));
    LocalMux I__1450 (
            .O(N__10524),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__1449 (
            .O(N__10519),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__1448 (
            .O(N__10514),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__1447 (
            .O(N__10511),
            .I(N__10506));
    InMux I__1446 (
            .O(N__10510),
            .I(N__10501));
    InMux I__1445 (
            .O(N__10509),
            .I(N__10501));
    LocalMux I__1444 (
            .O(N__10506),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__1443 (
            .O(N__10501),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__1442 (
            .O(N__10496),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__1441 (
            .O(N__10493),
            .I(\delay_measurement_inst.delay_hc_timer.N_105_cascade_ ));
    InMux I__1440 (
            .O(N__10490),
            .I(N__10485));
    InMux I__1439 (
            .O(N__10489),
            .I(N__10482));
    InMux I__1438 (
            .O(N__10488),
            .I(N__10479));
    LocalMux I__1437 (
            .O(N__10485),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__1436 (
            .O(N__10482),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__1435 (
            .O(N__10479),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__1434 (
            .O(N__10472),
            .I(N__10467));
    InMux I__1433 (
            .O(N__10471),
            .I(N__10464));
    InMux I__1432 (
            .O(N__10470),
            .I(N__10461));
    LocalMux I__1431 (
            .O(N__10467),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__1430 (
            .O(N__10464),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__1429 (
            .O(N__10461),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__1428 (
            .O(N__10454),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__1427 (
            .O(N__10451),
            .I(N__10446));
    CascadeMux I__1426 (
            .O(N__10450),
            .I(N__10443));
    InMux I__1425 (
            .O(N__10449),
            .I(N__10440));
    InMux I__1424 (
            .O(N__10446),
            .I(N__10435));
    InMux I__1423 (
            .O(N__10443),
            .I(N__10435));
    LocalMux I__1422 (
            .O(N__10440),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__1421 (
            .O(N__10435),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__1420 (
            .O(N__10430),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__1419 (
            .O(N__10427),
            .I(N__10422));
    CascadeMux I__1418 (
            .O(N__10426),
            .I(N__10419));
    InMux I__1417 (
            .O(N__10425),
            .I(N__10416));
    InMux I__1416 (
            .O(N__10422),
            .I(N__10411));
    InMux I__1415 (
            .O(N__10419),
            .I(N__10411));
    LocalMux I__1414 (
            .O(N__10416),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__1413 (
            .O(N__10411),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__1412 (
            .O(N__10406),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__1411 (
            .O(N__10403),
            .I(N__10398));
    InMux I__1410 (
            .O(N__10402),
            .I(N__10393));
    InMux I__1409 (
            .O(N__10401),
            .I(N__10393));
    LocalMux I__1408 (
            .O(N__10398),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__1407 (
            .O(N__10393),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__1406 (
            .O(N__10388),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__1405 (
            .O(N__10385),
            .I(N__10382));
    LocalMux I__1404 (
            .O(N__10382),
            .I(N__10379));
    Odrv12 I__1403 (
            .O(N__10379),
            .I(il_max_comp1_c));
    InMux I__1402 (
            .O(N__10376),
            .I(N__10373));
    LocalMux I__1401 (
            .O(N__10373),
            .I(N__10370));
    Span4Mux_h I__1400 (
            .O(N__10370),
            .I(N__10367));
    Odrv4 I__1399 (
            .O(N__10367),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__1398 (
            .O(N__10364),
            .I(N__10361));
    InMux I__1397 (
            .O(N__10361),
            .I(N__10358));
    LocalMux I__1396 (
            .O(N__10358),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__1395 (
            .O(N__10355),
            .I(N__10352));
    InMux I__1394 (
            .O(N__10352),
            .I(N__10349));
    LocalMux I__1393 (
            .O(N__10349),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__1392 (
            .O(N__10346),
            .I(N__10343));
    InMux I__1391 (
            .O(N__10343),
            .I(N__10340));
    LocalMux I__1390 (
            .O(N__10340),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    InMux I__1389 (
            .O(N__10337),
            .I(N__10334));
    LocalMux I__1388 (
            .O(N__10334),
            .I(N__10331));
    Odrv4 I__1387 (
            .O(N__10331),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__1386 (
            .O(N__10328),
            .I(N__10325));
    InMux I__1385 (
            .O(N__10325),
            .I(N__10322));
    LocalMux I__1384 (
            .O(N__10322),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__1383 (
            .O(N__10319),
            .I(N__10316));
    LocalMux I__1382 (
            .O(N__10316),
            .I(N__10313));
    Span4Mux_h I__1381 (
            .O(N__10313),
            .I(N__10310));
    Odrv4 I__1380 (
            .O(N__10310),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__1379 (
            .O(N__10307),
            .I(N__10304));
    InMux I__1378 (
            .O(N__10304),
            .I(N__10301));
    LocalMux I__1377 (
            .O(N__10301),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__1376 (
            .O(N__10298),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__1375 (
            .O(N__10295),
            .I(N__10292));
    InMux I__1374 (
            .O(N__10292),
            .I(N__10289));
    LocalMux I__1373 (
            .O(N__10289),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__1372 (
            .O(N__10286),
            .I(N__10283));
    InMux I__1371 (
            .O(N__10283),
            .I(N__10280));
    LocalMux I__1370 (
            .O(N__10280),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__1369 (
            .O(N__10277),
            .I(N__10274));
    LocalMux I__1368 (
            .O(N__10274),
            .I(N__10271));
    Odrv12 I__1367 (
            .O(N__10271),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__1366 (
            .O(N__10268),
            .I(N__10265));
    InMux I__1365 (
            .O(N__10265),
            .I(N__10262));
    LocalMux I__1364 (
            .O(N__10262),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__1363 (
            .O(N__10259),
            .I(N__10256));
    LocalMux I__1362 (
            .O(N__10256),
            .I(N__10253));
    Span4Mux_h I__1361 (
            .O(N__10253),
            .I(N__10250));
    Odrv4 I__1360 (
            .O(N__10250),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__1359 (
            .O(N__10247),
            .I(N__10244));
    InMux I__1358 (
            .O(N__10244),
            .I(N__10241));
    LocalMux I__1357 (
            .O(N__10241),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__1356 (
            .O(N__10238),
            .I(N__10235));
    LocalMux I__1355 (
            .O(N__10235),
            .I(N__10232));
    Odrv12 I__1354 (
            .O(N__10232),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__1353 (
            .O(N__10229),
            .I(N__10226));
    InMux I__1352 (
            .O(N__10226),
            .I(N__10223));
    LocalMux I__1351 (
            .O(N__10223),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__1350 (
            .O(N__10220),
            .I(N__10217));
    LocalMux I__1349 (
            .O(N__10217),
            .I(N__10214));
    Span4Mux_h I__1348 (
            .O(N__10214),
            .I(N__10211));
    Odrv4 I__1347 (
            .O(N__10211),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__1346 (
            .O(N__10208),
            .I(N__10205));
    InMux I__1345 (
            .O(N__10205),
            .I(N__10202));
    LocalMux I__1344 (
            .O(N__10202),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__1343 (
            .O(N__10199),
            .I(N__10196));
    LocalMux I__1342 (
            .O(N__10196),
            .I(N__10193));
    Odrv4 I__1341 (
            .O(N__10193),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__1340 (
            .O(N__10190),
            .I(N__10187));
    InMux I__1339 (
            .O(N__10187),
            .I(N__10184));
    LocalMux I__1338 (
            .O(N__10184),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__1337 (
            .O(N__10181),
            .I(N__10178));
    LocalMux I__1336 (
            .O(N__10178),
            .I(N__10175));
    Span4Mux_v I__1335 (
            .O(N__10175),
            .I(N__10172));
    Odrv4 I__1334 (
            .O(N__10172),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__1333 (
            .O(N__10169),
            .I(N__10166));
    InMux I__1332 (
            .O(N__10166),
            .I(N__10163));
    LocalMux I__1331 (
            .O(N__10163),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__1330 (
            .O(N__10160),
            .I(N__10152));
    InMux I__1329 (
            .O(N__10159),
            .I(N__10152));
    InMux I__1328 (
            .O(N__10158),
            .I(N__10147));
    InMux I__1327 (
            .O(N__10157),
            .I(N__10147));
    LocalMux I__1326 (
            .O(N__10152),
            .I(N__10144));
    LocalMux I__1325 (
            .O(N__10147),
            .I(N__10141));
    Odrv4 I__1324 (
            .O(N__10144),
            .I(\phase_controller_inst1.stoper_tr.un1_start ));
    Odrv4 I__1323 (
            .O(N__10141),
            .I(\phase_controller_inst1.stoper_tr.un1_start ));
    InMux I__1322 (
            .O(N__10136),
            .I(N__10133));
    LocalMux I__1321 (
            .O(N__10133),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__1320 (
            .O(N__10130),
            .I(N__10127));
    InMux I__1319 (
            .O(N__10127),
            .I(N__10124));
    LocalMux I__1318 (
            .O(N__10124),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__1317 (
            .O(N__10121),
            .I(N__10118));
    LocalMux I__1316 (
            .O(N__10118),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__1315 (
            .O(N__10115),
            .I(N__10112));
    InMux I__1314 (
            .O(N__10112),
            .I(N__10109));
    LocalMux I__1313 (
            .O(N__10109),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__1312 (
            .O(N__10106),
            .I(N__10103));
    LocalMux I__1311 (
            .O(N__10103),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__1310 (
            .O(N__10100),
            .I(N__10097));
    InMux I__1309 (
            .O(N__10097),
            .I(N__10094));
    LocalMux I__1308 (
            .O(N__10094),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__1307 (
            .O(N__10091),
            .I(N__10088));
    InMux I__1306 (
            .O(N__10088),
            .I(N__10085));
    LocalMux I__1305 (
            .O(N__10085),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__1304 (
            .O(N__10082),
            .I(N__10079));
    LocalMux I__1303 (
            .O(N__10079),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__1302 (
            .O(N__10076),
            .I(N__10073));
    InMux I__1301 (
            .O(N__10073),
            .I(N__10070));
    LocalMux I__1300 (
            .O(N__10070),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__1299 (
            .O(N__10067),
            .I(N__10064));
    LocalMux I__1298 (
            .O(N__10064),
            .I(N__10061));
    Odrv4 I__1297 (
            .O(N__10061),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ1Z_6 ));
    CascadeMux I__1296 (
            .O(N__10058),
            .I(N__10055));
    InMux I__1295 (
            .O(N__10055),
            .I(N__10052));
    LocalMux I__1294 (
            .O(N__10052),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__1293 (
            .O(N__10049),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto6Z0Z_0_cascade_ ));
    InMux I__1292 (
            .O(N__10046),
            .I(N__10043));
    LocalMux I__1291 (
            .O(N__10043),
            .I(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_4 ));
    CascadeMux I__1290 (
            .O(N__10040),
            .I(\phase_controller_inst1.stoper_tr.un2_startlt19_0_cascade_ ));
    InMux I__1289 (
            .O(N__10037),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__1288 (
            .O(N__10034),
            .I(bfn_7_19_0_));
    InMux I__1287 (
            .O(N__10031),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__1286 (
            .O(N__10028),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ));
    CascadeMux I__1285 (
            .O(N__10025),
            .I(\phase_controller_inst1.stoper_tr.un1_startlt8_cascade_ ));
    InMux I__1284 (
            .O(N__10022),
            .I(N__10019));
    LocalMux I__1283 (
            .O(N__10019),
            .I(\phase_controller_inst1.stoper_tr.un1_startlto5Z0Z_1 ));
    InMux I__1282 (
            .O(N__10016),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__1281 (
            .O(N__10013),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__1280 (
            .O(N__10010),
            .I(bfn_7_18_0_));
    InMux I__1279 (
            .O(N__10007),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__1278 (
            .O(N__10004),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__1277 (
            .O(N__10001),
            .I(N__9998));
    LocalMux I__1276 (
            .O(N__9998),
            .I(N__9995));
    Odrv4 I__1275 (
            .O(N__9995),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__1274 (
            .O(N__9992),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__1273 (
            .O(N__9989),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__1272 (
            .O(N__9986),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__1271 (
            .O(N__9983),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__1270 (
            .O(N__9980),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__1269 (
            .O(N__9977),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__1268 (
            .O(N__9974),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__1267 (
            .O(N__9971),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__1266 (
            .O(N__9968),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__1265 (
            .O(N__9965),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__1264 (
            .O(N__9962),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__1263 (
            .O(N__9959),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__1262 (
            .O(N__9956),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__1261 (
            .O(N__9953),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__1260 (
            .O(N__9950),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__1259 (
            .O(N__9947),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__1258 (
            .O(N__9944),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__1257 (
            .O(N__9941),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__1256 (
            .O(N__9938),
            .I(bfn_7_16_0_));
    InMux I__1255 (
            .O(N__9935),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__1254 (
            .O(N__9932),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__1253 (
            .O(N__9929),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__1252 (
            .O(N__9926),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__1251 (
            .O(N__9923),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__1250 (
            .O(N__9920),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__1249 (
            .O(N__9917),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__1248 (
            .O(N__9914),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__1247 (
            .O(N__9911),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__1246 (
            .O(N__9908),
            .I(bfn_7_15_0_));
    InMux I__1245 (
            .O(N__9905),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__1244 (
            .O(N__9902),
            .I(bfn_7_13_0_));
    InMux I__1243 (
            .O(N__9899),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__1242 (
            .O(N__9896),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__1241 (
            .O(N__9893),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__1240 (
            .O(N__9890),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__1239 (
            .O(N__9887),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__1238 (
            .O(N__9884),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__1237 (
            .O(N__9881),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__1236 (
            .O(N__9878),
            .I(bfn_7_14_0_));
    CascadeMux I__1235 (
            .O(N__9875),
            .I(N__9872));
    InMux I__1234 (
            .O(N__9872),
            .I(N__9869));
    LocalMux I__1233 (
            .O(N__9869),
            .I(\phase_controller_slave.stoper_hc.N_60 ));
    InMux I__1232 (
            .O(N__9866),
            .I(N__9858));
    InMux I__1231 (
            .O(N__9865),
            .I(N__9858));
    InMux I__1230 (
            .O(N__9864),
            .I(N__9855));
    InMux I__1229 (
            .O(N__9863),
            .I(N__9852));
    LocalMux I__1228 (
            .O(N__9858),
            .I(N__9847));
    LocalMux I__1227 (
            .O(N__9855),
            .I(N__9847));
    LocalMux I__1226 (
            .O(N__9852),
            .I(\phase_controller_slave.hc_time_passed ));
    Odrv4 I__1225 (
            .O(N__9847),
            .I(\phase_controller_slave.hc_time_passed ));
    InMux I__1224 (
            .O(N__9842),
            .I(N__9839));
    LocalMux I__1223 (
            .O(N__9839),
            .I(N__9835));
    InMux I__1222 (
            .O(N__9838),
            .I(N__9832));
    Odrv4 I__1221 (
            .O(N__9835),
            .I(\phase_controller_slave.state_RNIVDE2Z0Z_0 ));
    LocalMux I__1220 (
            .O(N__9832),
            .I(\phase_controller_slave.state_RNIVDE2Z0Z_0 ));
    CascadeMux I__1219 (
            .O(N__9827),
            .I(N__9824));
    InMux I__1218 (
            .O(N__9824),
            .I(N__9819));
    CascadeMux I__1217 (
            .O(N__9823),
            .I(N__9816));
    CascadeMux I__1216 (
            .O(N__9822),
            .I(N__9813));
    LocalMux I__1215 (
            .O(N__9819),
            .I(N__9809));
    InMux I__1214 (
            .O(N__9816),
            .I(N__9806));
    InMux I__1213 (
            .O(N__9813),
            .I(N__9801));
    InMux I__1212 (
            .O(N__9812),
            .I(N__9801));
    Span4Mux_h I__1211 (
            .O(N__9809),
            .I(N__9798));
    LocalMux I__1210 (
            .O(N__9806),
            .I(N__9795));
    LocalMux I__1209 (
            .O(N__9801),
            .I(N__9792));
    Odrv4 I__1208 (
            .O(N__9798),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    Odrv4 I__1207 (
            .O(N__9795),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    Odrv4 I__1206 (
            .O(N__9792),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    InMux I__1205 (
            .O(N__9785),
            .I(N__9782));
    LocalMux I__1204 (
            .O(N__9782),
            .I(\phase_controller_slave.state_RNO_0Z0Z_3 ));
    InMux I__1203 (
            .O(N__9779),
            .I(N__9775));
    CascadeMux I__1202 (
            .O(N__9778),
            .I(N__9772));
    LocalMux I__1201 (
            .O(N__9775),
            .I(N__9768));
    InMux I__1200 (
            .O(N__9772),
            .I(N__9765));
    InMux I__1199 (
            .O(N__9771),
            .I(N__9762));
    Odrv4 I__1198 (
            .O(N__9768),
            .I(shift_flag_start));
    LocalMux I__1197 (
            .O(N__9765),
            .I(shift_flag_start));
    LocalMux I__1196 (
            .O(N__9762),
            .I(shift_flag_start));
    InMux I__1195 (
            .O(N__9755),
            .I(N__9752));
    LocalMux I__1194 (
            .O(N__9752),
            .I(N__9746));
    InMux I__1193 (
            .O(N__9751),
            .I(N__9743));
    InMux I__1192 (
            .O(N__9750),
            .I(N__9740));
    InMux I__1191 (
            .O(N__9749),
            .I(N__9737));
    Odrv12 I__1190 (
            .O(N__9746),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    LocalMux I__1189 (
            .O(N__9743),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    LocalMux I__1188 (
            .O(N__9740),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    LocalMux I__1187 (
            .O(N__9737),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    IoInMux I__1186 (
            .O(N__9728),
            .I(N__9725));
    LocalMux I__1185 (
            .O(N__9725),
            .I(N__9722));
    IoSpan4Mux I__1184 (
            .O(N__9722),
            .I(N__9719));
    Span4Mux_s2_v I__1183 (
            .O(N__9719),
            .I(N__9716));
    Span4Mux_v I__1182 (
            .O(N__9716),
            .I(N__9713));
    Odrv4 I__1181 (
            .O(N__9713),
            .I(s4_phy_c));
    InMux I__1180 (
            .O(N__9710),
            .I(N__9707));
    LocalMux I__1179 (
            .O(N__9707),
            .I(N__9704));
    Odrv4 I__1178 (
            .O(N__9704),
            .I(il_max_comp2_D1));
    InMux I__1177 (
            .O(N__9701),
            .I(N__9698));
    LocalMux I__1176 (
            .O(N__9698),
            .I(N__9695));
    Odrv4 I__1175 (
            .O(N__9695),
            .I(\phase_controller_slave.start_timer_hc_0_sqmuxa ));
    InMux I__1174 (
            .O(N__9692),
            .I(N__9689));
    LocalMux I__1173 (
            .O(N__9689),
            .I(\phase_controller_slave.start_timer_hc_RNOZ0Z_0 ));
    InMux I__1172 (
            .O(N__9686),
            .I(N__9681));
    InMux I__1171 (
            .O(N__9685),
            .I(N__9678));
    InMux I__1170 (
            .O(N__9684),
            .I(N__9675));
    LocalMux I__1169 (
            .O(N__9681),
            .I(N__9668));
    LocalMux I__1168 (
            .O(N__9678),
            .I(N__9668));
    LocalMux I__1167 (
            .O(N__9675),
            .I(N__9668));
    Span4Mux_v I__1166 (
            .O(N__9668),
            .I(N__9665));
    Odrv4 I__1165 (
            .O(N__9665),
            .I(il_min_comp2_D2));
    CascadeMux I__1164 (
            .O(N__9662),
            .I(N__9659));
    InMux I__1163 (
            .O(N__9659),
            .I(N__9652));
    InMux I__1162 (
            .O(N__9658),
            .I(N__9652));
    InMux I__1161 (
            .O(N__9657),
            .I(N__9649));
    LocalMux I__1160 (
            .O(N__9652),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    LocalMux I__1159 (
            .O(N__9649),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    InMux I__1158 (
            .O(N__9644),
            .I(N__9640));
    InMux I__1157 (
            .O(N__9643),
            .I(N__9637));
    LocalMux I__1156 (
            .O(N__9640),
            .I(N__9631));
    LocalMux I__1155 (
            .O(N__9637),
            .I(N__9631));
    InMux I__1154 (
            .O(N__9636),
            .I(N__9628));
    Odrv12 I__1153 (
            .O(N__9631),
            .I(il_max_comp2_D2));
    LocalMux I__1152 (
            .O(N__9628),
            .I(il_max_comp2_D2));
    InMux I__1151 (
            .O(N__9623),
            .I(N__9620));
    LocalMux I__1150 (
            .O(N__9620),
            .I(N__9617));
    Odrv4 I__1149 (
            .O(N__9617),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ));
    InMux I__1148 (
            .O(N__9614),
            .I(N__9611));
    LocalMux I__1147 (
            .O(N__9611),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ));
    InMux I__1146 (
            .O(N__9608),
            .I(N__9605));
    LocalMux I__1145 (
            .O(N__9605),
            .I(N__9602));
    Odrv4 I__1144 (
            .O(N__9602),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ));
    InMux I__1143 (
            .O(N__9599),
            .I(N__9596));
    LocalMux I__1142 (
            .O(N__9596),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ));
    InMux I__1141 (
            .O(N__9593),
            .I(N__9590));
    LocalMux I__1140 (
            .O(N__9590),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ));
    CEMux I__1139 (
            .O(N__9587),
            .I(N__9584));
    LocalMux I__1138 (
            .O(N__9584),
            .I(N__9579));
    CEMux I__1137 (
            .O(N__9583),
            .I(N__9576));
    CEMux I__1136 (
            .O(N__9582),
            .I(N__9572));
    Span4Mux_h I__1135 (
            .O(N__9579),
            .I(N__9567));
    LocalMux I__1134 (
            .O(N__9576),
            .I(N__9567));
    CEMux I__1133 (
            .O(N__9575),
            .I(N__9564));
    LocalMux I__1132 (
            .O(N__9572),
            .I(N__9561));
    Span4Mux_v I__1131 (
            .O(N__9567),
            .I(N__9558));
    LocalMux I__1130 (
            .O(N__9564),
            .I(N__9555));
    Span4Mux_h I__1129 (
            .O(N__9561),
            .I(N__9552));
    Span4Mux_h I__1128 (
            .O(N__9558),
            .I(N__9549));
    Span4Mux_h I__1127 (
            .O(N__9555),
            .I(N__9546));
    Odrv4 I__1126 (
            .O(N__9552),
            .I(\phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1 ));
    Odrv4 I__1125 (
            .O(N__9549),
            .I(\phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1 ));
    Odrv4 I__1124 (
            .O(N__9546),
            .I(\phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1 ));
    InMux I__1123 (
            .O(N__9539),
            .I(N__9536));
    LocalMux I__1122 (
            .O(N__9536),
            .I(N__9533));
    Span12Mux_v I__1121 (
            .O(N__9533),
            .I(N__9530));
    Odrv12 I__1120 (
            .O(N__9530),
            .I(il_max_comp2_c));
    InMux I__1119 (
            .O(N__9527),
            .I(N__9524));
    LocalMux I__1118 (
            .O(N__9524),
            .I(N__9521));
    Span4Mux_h I__1117 (
            .O(N__9521),
            .I(N__9518));
    Span4Mux_v I__1116 (
            .O(N__9518),
            .I(N__9515));
    Span4Mux_v I__1115 (
            .O(N__9515),
            .I(N__9512));
    Odrv4 I__1114 (
            .O(N__9512),
            .I(il_min_comp2_c));
    InMux I__1113 (
            .O(N__9509),
            .I(N__9506));
    LocalMux I__1112 (
            .O(N__9506),
            .I(il_min_comp2_D1));
    InMux I__1111 (
            .O(N__9503),
            .I(N__9500));
    LocalMux I__1110 (
            .O(N__9500),
            .I(N__9497));
    Odrv4 I__1109 (
            .O(N__9497),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ));
    InMux I__1108 (
            .O(N__9494),
            .I(N__9491));
    LocalMux I__1107 (
            .O(N__9491),
            .I(N__9488));
    Odrv4 I__1106 (
            .O(N__9488),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ));
    InMux I__1105 (
            .O(N__9485),
            .I(N__9482));
    LocalMux I__1104 (
            .O(N__9482),
            .I(N__9479));
    Odrv4 I__1103 (
            .O(N__9479),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ));
    InMux I__1102 (
            .O(N__9476),
            .I(N__9473));
    LocalMux I__1101 (
            .O(N__9473),
            .I(N__9470));
    Span4Mux_h I__1100 (
            .O(N__9470),
            .I(N__9467));
    Odrv4 I__1099 (
            .O(N__9467),
            .I(\phase_controller_slave.stoper_tr.target_timeZ1Z_6 ));
    InMux I__1098 (
            .O(N__9464),
            .I(N__9461));
    LocalMux I__1097 (
            .O(N__9461),
            .I(N__9458));
    Odrv4 I__1096 (
            .O(N__9458),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ));
    InMux I__1095 (
            .O(N__9455),
            .I(N__9452));
    LocalMux I__1094 (
            .O(N__9452),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ));
    InMux I__1093 (
            .O(N__9449),
            .I(N__9446));
    LocalMux I__1092 (
            .O(N__9446),
            .I(N__9443));
    Span4Mux_v I__1091 (
            .O(N__9443),
            .I(N__9440));
    Odrv4 I__1090 (
            .O(N__9440),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ));
    InMux I__1089 (
            .O(N__9437),
            .I(N__9434));
    LocalMux I__1088 (
            .O(N__9434),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ));
    InMux I__1087 (
            .O(N__9431),
            .I(N__9428));
    LocalMux I__1086 (
            .O(N__9428),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ));
    InMux I__1085 (
            .O(N__9425),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__1084 (
            .O(N__9422),
            .I(N__9419));
    LocalMux I__1083 (
            .O(N__9419),
            .I(N__9411));
    InMux I__1082 (
            .O(N__9418),
            .I(N__9400));
    InMux I__1081 (
            .O(N__9417),
            .I(N__9400));
    InMux I__1080 (
            .O(N__9416),
            .I(N__9400));
    InMux I__1079 (
            .O(N__9415),
            .I(N__9400));
    InMux I__1078 (
            .O(N__9414),
            .I(N__9400));
    Odrv4 I__1077 (
            .O(N__9411),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__1076 (
            .O(N__9400),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__1075 (
            .O(N__9395),
            .I(N__9392));
    InMux I__1074 (
            .O(N__9392),
            .I(N__9387));
    InMux I__1073 (
            .O(N__9391),
            .I(N__9384));
    InMux I__1072 (
            .O(N__9390),
            .I(N__9381));
    LocalMux I__1071 (
            .O(N__9387),
            .I(\phase_controller_slave.tr_time_passed ));
    LocalMux I__1070 (
            .O(N__9384),
            .I(\phase_controller_slave.tr_time_passed ));
    LocalMux I__1069 (
            .O(N__9381),
            .I(\phase_controller_slave.tr_time_passed ));
    InMux I__1068 (
            .O(N__9374),
            .I(N__9370));
    InMux I__1067 (
            .O(N__9373),
            .I(N__9367));
    LocalMux I__1066 (
            .O(N__9370),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    LocalMux I__1065 (
            .O(N__9367),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    InMux I__1064 (
            .O(N__9362),
            .I(N__9359));
    LocalMux I__1063 (
            .O(N__9359),
            .I(\phase_controller_slave.start_timer_tr_0_sqmuxa ));
    InMux I__1062 (
            .O(N__9356),
            .I(N__9353));
    LocalMux I__1061 (
            .O(N__9353),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ));
    InMux I__1060 (
            .O(N__9350),
            .I(N__9347));
    LocalMux I__1059 (
            .O(N__9347),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ));
    InMux I__1058 (
            .O(N__9344),
            .I(N__9341));
    LocalMux I__1057 (
            .O(N__9341),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ));
    InMux I__1056 (
            .O(N__9338),
            .I(N__9335));
    LocalMux I__1055 (
            .O(N__9335),
            .I(N__9332));
    Odrv4 I__1054 (
            .O(N__9332),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ));
    InMux I__1053 (
            .O(N__9329),
            .I(N__9326));
    LocalMux I__1052 (
            .O(N__9326),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ));
    InMux I__1051 (
            .O(N__9323),
            .I(N__9319));
    InMux I__1050 (
            .O(N__9322),
            .I(N__9316));
    LocalMux I__1049 (
            .O(N__9319),
            .I(N__9313));
    LocalMux I__1048 (
            .O(N__9316),
            .I(N__9310));
    Span4Mux_v I__1047 (
            .O(N__9313),
            .I(N__9307));
    Span4Mux_v I__1046 (
            .O(N__9310),
            .I(N__9304));
    Odrv4 I__1045 (
            .O(N__9307),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__1044 (
            .O(N__9304),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__1043 (
            .O(N__9299),
            .I(N__9296));
    InMux I__1042 (
            .O(N__9296),
            .I(N__9293));
    LocalMux I__1041 (
            .O(N__9293),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ));
    InMux I__1040 (
            .O(N__9290),
            .I(N__9286));
    InMux I__1039 (
            .O(N__9289),
            .I(N__9283));
    LocalMux I__1038 (
            .O(N__9286),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__1037 (
            .O(N__9283),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__1036 (
            .O(N__9278),
            .I(N__9275));
    InMux I__1035 (
            .O(N__9275),
            .I(N__9272));
    LocalMux I__1034 (
            .O(N__9272),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ));
    InMux I__1033 (
            .O(N__9269),
            .I(N__9265));
    InMux I__1032 (
            .O(N__9268),
            .I(N__9262));
    LocalMux I__1031 (
            .O(N__9265),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__1030 (
            .O(N__9262),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__1029 (
            .O(N__9257),
            .I(N__9254));
    InMux I__1028 (
            .O(N__9254),
            .I(N__9251));
    LocalMux I__1027 (
            .O(N__9251),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ));
    InMux I__1026 (
            .O(N__9248),
            .I(N__9244));
    InMux I__1025 (
            .O(N__9247),
            .I(N__9241));
    LocalMux I__1024 (
            .O(N__9244),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__1023 (
            .O(N__9241),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__1022 (
            .O(N__9236),
            .I(N__9233));
    InMux I__1021 (
            .O(N__9233),
            .I(N__9230));
    LocalMux I__1020 (
            .O(N__9230),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ));
    InMux I__1019 (
            .O(N__9227),
            .I(N__9223));
    InMux I__1018 (
            .O(N__9226),
            .I(N__9220));
    LocalMux I__1017 (
            .O(N__9223),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__1016 (
            .O(N__9220),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__1015 (
            .O(N__9215),
            .I(N__9212));
    InMux I__1014 (
            .O(N__9212),
            .I(N__9209));
    LocalMux I__1013 (
            .O(N__9209),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ));
    InMux I__1012 (
            .O(N__9206),
            .I(N__9202));
    InMux I__1011 (
            .O(N__9205),
            .I(N__9199));
    LocalMux I__1010 (
            .O(N__9202),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__1009 (
            .O(N__9199),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__1008 (
            .O(N__9194),
            .I(N__9191));
    InMux I__1007 (
            .O(N__9191),
            .I(N__9188));
    LocalMux I__1006 (
            .O(N__9188),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ));
    InMux I__1005 (
            .O(N__9185),
            .I(N__9181));
    InMux I__1004 (
            .O(N__9184),
            .I(N__9178));
    LocalMux I__1003 (
            .O(N__9181),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__1002 (
            .O(N__9178),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    CascadeMux I__1001 (
            .O(N__9173),
            .I(N__9170));
    InMux I__1000 (
            .O(N__9170),
            .I(N__9167));
    LocalMux I__999 (
            .O(N__9167),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ));
    InMux I__998 (
            .O(N__9164),
            .I(N__9160));
    InMux I__997 (
            .O(N__9163),
            .I(N__9157));
    LocalMux I__996 (
            .O(N__9160),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__995 (
            .O(N__9157),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__994 (
            .O(N__9152),
            .I(N__9149));
    InMux I__993 (
            .O(N__9149),
            .I(N__9146));
    LocalMux I__992 (
            .O(N__9146),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ));
    InMux I__991 (
            .O(N__9143),
            .I(N__9139));
    InMux I__990 (
            .O(N__9142),
            .I(N__9136));
    LocalMux I__989 (
            .O(N__9139),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__988 (
            .O(N__9136),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__987 (
            .O(N__9131),
            .I(N__9128));
    InMux I__986 (
            .O(N__9128),
            .I(N__9125));
    LocalMux I__985 (
            .O(N__9125),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ));
    InMux I__984 (
            .O(N__9122),
            .I(N__9119));
    LocalMux I__983 (
            .O(N__9119),
            .I(N__9115));
    InMux I__982 (
            .O(N__9118),
            .I(N__9112));
    Odrv4 I__981 (
            .O(N__9115),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__980 (
            .O(N__9112),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__979 (
            .O(N__9107),
            .I(N__9104));
    InMux I__978 (
            .O(N__9104),
            .I(N__9101));
    LocalMux I__977 (
            .O(N__9101),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__976 (
            .O(N__9098),
            .I(N__9095));
    InMux I__975 (
            .O(N__9095),
            .I(N__9091));
    InMux I__974 (
            .O(N__9094),
            .I(N__9088));
    LocalMux I__973 (
            .O(N__9091),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__972 (
            .O(N__9088),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__971 (
            .O(N__9083),
            .I(N__9080));
    InMux I__970 (
            .O(N__9080),
            .I(N__9077));
    LocalMux I__969 (
            .O(N__9077),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ));
    InMux I__968 (
            .O(N__9074),
            .I(N__9070));
    InMux I__967 (
            .O(N__9073),
            .I(N__9067));
    LocalMux I__966 (
            .O(N__9070),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__965 (
            .O(N__9067),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__964 (
            .O(N__9062),
            .I(N__9059));
    InMux I__963 (
            .O(N__9059),
            .I(N__9056));
    LocalMux I__962 (
            .O(N__9056),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__961 (
            .O(N__9053),
            .I(N__9050));
    InMux I__960 (
            .O(N__9050),
            .I(N__9046));
    InMux I__959 (
            .O(N__9049),
            .I(N__9043));
    LocalMux I__958 (
            .O(N__9046),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__957 (
            .O(N__9043),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__956 (
            .O(N__9038),
            .I(N__9035));
    InMux I__955 (
            .O(N__9035),
            .I(N__9032));
    LocalMux I__954 (
            .O(N__9032),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ));
    InMux I__953 (
            .O(N__9029),
            .I(N__9025));
    InMux I__952 (
            .O(N__9028),
            .I(N__9022));
    LocalMux I__951 (
            .O(N__9025),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__950 (
            .O(N__9022),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__949 (
            .O(N__9017),
            .I(N__9014));
    InMux I__948 (
            .O(N__9014),
            .I(N__9011));
    LocalMux I__947 (
            .O(N__9011),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ));
    InMux I__946 (
            .O(N__9008),
            .I(N__9004));
    InMux I__945 (
            .O(N__9007),
            .I(N__9001));
    LocalMux I__944 (
            .O(N__9004),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__943 (
            .O(N__9001),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__942 (
            .O(N__8996),
            .I(N__8993));
    InMux I__941 (
            .O(N__8993),
            .I(N__8990));
    LocalMux I__940 (
            .O(N__8990),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ));
    InMux I__939 (
            .O(N__8987),
            .I(N__8983));
    InMux I__938 (
            .O(N__8986),
            .I(N__8980));
    LocalMux I__937 (
            .O(N__8983),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__936 (
            .O(N__8980),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    CascadeMux I__935 (
            .O(N__8975),
            .I(N__8972));
    InMux I__934 (
            .O(N__8972),
            .I(N__8969));
    LocalMux I__933 (
            .O(N__8969),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ));
    InMux I__932 (
            .O(N__8966),
            .I(N__8963));
    LocalMux I__931 (
            .O(N__8963),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ));
    InMux I__930 (
            .O(N__8960),
            .I(N__8957));
    LocalMux I__929 (
            .O(N__8957),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ));
    CascadeMux I__928 (
            .O(N__8954),
            .I(N__8942));
    CascadeMux I__927 (
            .O(N__8953),
            .I(N__8935));
    CascadeMux I__926 (
            .O(N__8952),
            .I(N__8932));
    CascadeMux I__925 (
            .O(N__8951),
            .I(N__8929));
    CascadeMux I__924 (
            .O(N__8950),
            .I(N__8923));
    CascadeMux I__923 (
            .O(N__8949),
            .I(N__8920));
    CascadeMux I__922 (
            .O(N__8948),
            .I(N__8917));
    CascadeMux I__921 (
            .O(N__8947),
            .I(N__8914));
    CascadeMux I__920 (
            .O(N__8946),
            .I(N__8908));
    CascadeMux I__919 (
            .O(N__8945),
            .I(N__8905));
    InMux I__918 (
            .O(N__8942),
            .I(N__8899));
    InMux I__917 (
            .O(N__8941),
            .I(N__8884));
    InMux I__916 (
            .O(N__8940),
            .I(N__8884));
    InMux I__915 (
            .O(N__8939),
            .I(N__8884));
    InMux I__914 (
            .O(N__8938),
            .I(N__8884));
    InMux I__913 (
            .O(N__8935),
            .I(N__8884));
    InMux I__912 (
            .O(N__8932),
            .I(N__8884));
    InMux I__911 (
            .O(N__8929),
            .I(N__8884));
    InMux I__910 (
            .O(N__8928),
            .I(N__8881));
    InMux I__909 (
            .O(N__8927),
            .I(N__8876));
    InMux I__908 (
            .O(N__8926),
            .I(N__8876));
    InMux I__907 (
            .O(N__8923),
            .I(N__8861));
    InMux I__906 (
            .O(N__8920),
            .I(N__8861));
    InMux I__905 (
            .O(N__8917),
            .I(N__8861));
    InMux I__904 (
            .O(N__8914),
            .I(N__8861));
    InMux I__903 (
            .O(N__8913),
            .I(N__8861));
    InMux I__902 (
            .O(N__8912),
            .I(N__8861));
    InMux I__901 (
            .O(N__8911),
            .I(N__8861));
    InMux I__900 (
            .O(N__8908),
            .I(N__8850));
    InMux I__899 (
            .O(N__8905),
            .I(N__8850));
    InMux I__898 (
            .O(N__8904),
            .I(N__8850));
    InMux I__897 (
            .O(N__8903),
            .I(N__8850));
    InMux I__896 (
            .O(N__8902),
            .I(N__8850));
    LocalMux I__895 (
            .O(N__8899),
            .I(N__8847));
    LocalMux I__894 (
            .O(N__8884),
            .I(N__8840));
    LocalMux I__893 (
            .O(N__8881),
            .I(N__8840));
    LocalMux I__892 (
            .O(N__8876),
            .I(N__8840));
    LocalMux I__891 (
            .O(N__8861),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__890 (
            .O(N__8850),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__889 (
            .O(N__8847),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__888 (
            .O(N__8840),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__887 (
            .O(N__8831),
            .I(N__8828));
    LocalMux I__886 (
            .O(N__8828),
            .I(N__8825));
    Span4Mux_v I__885 (
            .O(N__8825),
            .I(N__8822));
    Odrv4 I__884 (
            .O(N__8822),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ));
    CascadeMux I__883 (
            .O(N__8819),
            .I(N__8813));
    CascadeMux I__882 (
            .O(N__8818),
            .I(N__8807));
    CascadeMux I__881 (
            .O(N__8817),
            .I(N__8804));
    CascadeMux I__880 (
            .O(N__8816),
            .I(N__8801));
    InMux I__879 (
            .O(N__8813),
            .I(N__8786));
    InMux I__878 (
            .O(N__8812),
            .I(N__8781));
    InMux I__877 (
            .O(N__8811),
            .I(N__8781));
    CascadeMux I__876 (
            .O(N__8810),
            .I(N__8774));
    InMux I__875 (
            .O(N__8807),
            .I(N__8766));
    InMux I__874 (
            .O(N__8804),
            .I(N__8766));
    InMux I__873 (
            .O(N__8801),
            .I(N__8766));
    InMux I__872 (
            .O(N__8800),
            .I(N__8763));
    InMux I__871 (
            .O(N__8799),
            .I(N__8746));
    InMux I__870 (
            .O(N__8798),
            .I(N__8746));
    InMux I__869 (
            .O(N__8797),
            .I(N__8746));
    InMux I__868 (
            .O(N__8796),
            .I(N__8746));
    InMux I__867 (
            .O(N__8795),
            .I(N__8746));
    InMux I__866 (
            .O(N__8794),
            .I(N__8746));
    InMux I__865 (
            .O(N__8793),
            .I(N__8746));
    InMux I__864 (
            .O(N__8792),
            .I(N__8737));
    InMux I__863 (
            .O(N__8791),
            .I(N__8737));
    InMux I__862 (
            .O(N__8790),
            .I(N__8737));
    InMux I__861 (
            .O(N__8789),
            .I(N__8737));
    LocalMux I__860 (
            .O(N__8786),
            .I(N__8734));
    LocalMux I__859 (
            .O(N__8781),
            .I(N__8731));
    InMux I__858 (
            .O(N__8780),
            .I(N__8718));
    InMux I__857 (
            .O(N__8779),
            .I(N__8718));
    InMux I__856 (
            .O(N__8778),
            .I(N__8718));
    InMux I__855 (
            .O(N__8777),
            .I(N__8718));
    InMux I__854 (
            .O(N__8774),
            .I(N__8718));
    InMux I__853 (
            .O(N__8773),
            .I(N__8718));
    LocalMux I__852 (
            .O(N__8766),
            .I(N__8713));
    LocalMux I__851 (
            .O(N__8763),
            .I(N__8713));
    InMux I__850 (
            .O(N__8762),
            .I(N__8708));
    InMux I__849 (
            .O(N__8761),
            .I(N__8708));
    LocalMux I__848 (
            .O(N__8746),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__847 (
            .O(N__8737),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__846 (
            .O(N__8734),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__845 (
            .O(N__8731),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__844 (
            .O(N__8718),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__843 (
            .O(N__8713),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__842 (
            .O(N__8708),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__841 (
            .O(N__8693),
            .I(N__8690));
    InMux I__840 (
            .O(N__8690),
            .I(N__8687));
    LocalMux I__839 (
            .O(N__8687),
            .I(\phase_controller_slave.stoper_tr.N_60 ));
    InMux I__838 (
            .O(N__8684),
            .I(N__8650));
    InMux I__837 (
            .O(N__8683),
            .I(N__8650));
    InMux I__836 (
            .O(N__8682),
            .I(N__8650));
    InMux I__835 (
            .O(N__8681),
            .I(N__8650));
    InMux I__834 (
            .O(N__8680),
            .I(N__8650));
    InMux I__833 (
            .O(N__8679),
            .I(N__8650));
    InMux I__832 (
            .O(N__8678),
            .I(N__8650));
    InMux I__831 (
            .O(N__8677),
            .I(N__8633));
    InMux I__830 (
            .O(N__8676),
            .I(N__8633));
    InMux I__829 (
            .O(N__8675),
            .I(N__8633));
    InMux I__828 (
            .O(N__8674),
            .I(N__8633));
    InMux I__827 (
            .O(N__8673),
            .I(N__8633));
    InMux I__826 (
            .O(N__8672),
            .I(N__8633));
    InMux I__825 (
            .O(N__8671),
            .I(N__8633));
    InMux I__824 (
            .O(N__8670),
            .I(N__8622));
    InMux I__823 (
            .O(N__8669),
            .I(N__8622));
    InMux I__822 (
            .O(N__8668),
            .I(N__8622));
    InMux I__821 (
            .O(N__8667),
            .I(N__8622));
    InMux I__820 (
            .O(N__8666),
            .I(N__8622));
    InMux I__819 (
            .O(N__8665),
            .I(N__8617));
    LocalMux I__818 (
            .O(N__8650),
            .I(N__8614));
    InMux I__817 (
            .O(N__8649),
            .I(N__8611));
    InMux I__816 (
            .O(N__8648),
            .I(N__8608));
    LocalMux I__815 (
            .O(N__8633),
            .I(N__8603));
    LocalMux I__814 (
            .O(N__8622),
            .I(N__8603));
    InMux I__813 (
            .O(N__8621),
            .I(N__8598));
    InMux I__812 (
            .O(N__8620),
            .I(N__8598));
    LocalMux I__811 (
            .O(N__8617),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__810 (
            .O(N__8614),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    LocalMux I__809 (
            .O(N__8611),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    LocalMux I__808 (
            .O(N__8608),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__807 (
            .O(N__8603),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    LocalMux I__806 (
            .O(N__8598),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    InMux I__805 (
            .O(N__8585),
            .I(N__8580));
    InMux I__804 (
            .O(N__8584),
            .I(N__8577));
    InMux I__803 (
            .O(N__8583),
            .I(N__8574));
    LocalMux I__802 (
            .O(N__8580),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__801 (
            .O(N__8577),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__800 (
            .O(N__8574),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__799 (
            .O(N__8567),
            .I(N__8564));
    InMux I__798 (
            .O(N__8564),
            .I(N__8561));
    LocalMux I__797 (
            .O(N__8561),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ));
    InMux I__796 (
            .O(N__8558),
            .I(N__8555));
    LocalMux I__795 (
            .O(N__8555),
            .I(N__8552));
    Span4Mux_s3_h I__794 (
            .O(N__8552),
            .I(N__8548));
    InMux I__793 (
            .O(N__8551),
            .I(N__8545));
    Odrv4 I__792 (
            .O(N__8548),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__791 (
            .O(N__8545),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    CascadeMux I__790 (
            .O(N__8540),
            .I(N__8537));
    InMux I__789 (
            .O(N__8537),
            .I(N__8534));
    LocalMux I__788 (
            .O(N__8534),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ));
    InMux I__787 (
            .O(N__8531),
            .I(N__8527));
    InMux I__786 (
            .O(N__8530),
            .I(N__8524));
    LocalMux I__785 (
            .O(N__8527),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__784 (
            .O(N__8524),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__783 (
            .O(N__8519),
            .I(N__8516));
    InMux I__782 (
            .O(N__8516),
            .I(N__8513));
    LocalMux I__781 (
            .O(N__8513),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__780 (
            .O(N__8510),
            .I(N__8507));
    InMux I__779 (
            .O(N__8507),
            .I(N__8504));
    LocalMux I__778 (
            .O(N__8504),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    CascadeMux I__777 (
            .O(N__8501),
            .I(N__8498));
    InMux I__776 (
            .O(N__8498),
            .I(N__8495));
    LocalMux I__775 (
            .O(N__8495),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUSZ0Z53 ));
    CascadeMux I__774 (
            .O(N__8492),
            .I(N__8489));
    InMux I__773 (
            .O(N__8489),
            .I(N__8486));
    LocalMux I__772 (
            .O(N__8486),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ));
    InMux I__771 (
            .O(N__8483),
            .I(N__8480));
    LocalMux I__770 (
            .O(N__8480),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ));
    InMux I__769 (
            .O(N__8477),
            .I(N__8474));
    LocalMux I__768 (
            .O(N__8474),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ));
    InMux I__767 (
            .O(N__8471),
            .I(N__8468));
    LocalMux I__766 (
            .O(N__8468),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ));
    InMux I__765 (
            .O(N__8465),
            .I(N__8462));
    LocalMux I__764 (
            .O(N__8462),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ));
    InMux I__763 (
            .O(N__8459),
            .I(N__8456));
    LocalMux I__762 (
            .O(N__8456),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__761 (
            .O(N__8453),
            .I(N__8450));
    LocalMux I__760 (
            .O(N__8450),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ));
    InMux I__759 (
            .O(N__8447),
            .I(N__8444));
    LocalMux I__758 (
            .O(N__8444),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ));
    CascadeMux I__757 (
            .O(N__8441),
            .I(N__8438));
    InMux I__756 (
            .O(N__8438),
            .I(N__8435));
    LocalMux I__755 (
            .O(N__8435),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ));
    InMux I__754 (
            .O(N__8432),
            .I(N__8429));
    LocalMux I__753 (
            .O(N__8429),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ));
    CascadeMux I__752 (
            .O(N__8426),
            .I(N__8423));
    InMux I__751 (
            .O(N__8423),
            .I(N__8420));
    LocalMux I__750 (
            .O(N__8420),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ));
    InMux I__749 (
            .O(N__8417),
            .I(N__8414));
    LocalMux I__748 (
            .O(N__8414),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ));
    CascadeMux I__747 (
            .O(N__8411),
            .I(N__8408));
    InMux I__746 (
            .O(N__8408),
            .I(N__8405));
    LocalMux I__745 (
            .O(N__8405),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ));
    CascadeMux I__744 (
            .O(N__8402),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    InMux I__743 (
            .O(N__8399),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__742 (
            .O(N__8396),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__741 (
            .O(N__8393),
            .I(N__8390));
    LocalMux I__740 (
            .O(N__8390),
            .I(N_39_i_i));
    InMux I__739 (
            .O(N__8387),
            .I(N__8384));
    LocalMux I__738 (
            .O(N__8384),
            .I(N__8381));
    Span12Mux_s3_v I__737 (
            .O(N__8381),
            .I(N__8378));
    Span12Mux_h I__736 (
            .O(N__8378),
            .I(N__8375));
    Span12Mux_h I__735 (
            .O(N__8375),
            .I(N__8369));
    InMux I__734 (
            .O(N__8374),
            .I(N__8366));
    InMux I__733 (
            .O(N__8373),
            .I(N__8363));
    InMux I__732 (
            .O(N__8372),
            .I(N__8360));
    Odrv12 I__731 (
            .O(N__8369),
            .I(CONSTANT_ONE_NET));
    LocalMux I__730 (
            .O(N__8366),
            .I(CONSTANT_ONE_NET));
    LocalMux I__729 (
            .O(N__8363),
            .I(CONSTANT_ONE_NET));
    LocalMux I__728 (
            .O(N__8360),
            .I(CONSTANT_ONE_NET));
    InMux I__727 (
            .O(N__8351),
            .I(N__8348));
    LocalMux I__726 (
            .O(N__8348),
            .I(rgb_drv_RNOZ0));
    InMux I__725 (
            .O(N__8345),
            .I(N__8342));
    LocalMux I__724 (
            .O(N__8342),
            .I(N__8339));
    Odrv4 I__723 (
            .O(N__8339),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ));
    CascadeMux I__722 (
            .O(N__8336),
            .I(N__8333));
    InMux I__721 (
            .O(N__8333),
            .I(N__8330));
    LocalMux I__720 (
            .O(N__8330),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ));
    InMux I__719 (
            .O(N__8327),
            .I(bfn_1_19_0_));
    InMux I__718 (
            .O(N__8324),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__717 (
            .O(N__8321),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__716 (
            .O(N__8318),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__715 (
            .O(N__8315),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__714 (
            .O(N__8312),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__713 (
            .O(N__8309),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__712 (
            .O(N__8306),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__711 (
            .O(N__8303),
            .I(bfn_1_20_0_));
    InMux I__710 (
            .O(N__8300),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__709 (
            .O(N__8297),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__708 (
            .O(N__8294),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__707 (
            .O(N__8291),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__706 (
            .O(N__8288),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__705 (
            .O(N__8285),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__704 (
            .O(N__8282),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_7_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_18_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_7_18_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_8_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_25_0_));
    defparam IN_MUX_bfv_8_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_26_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_8_26_0_));
    defparam IN_MUX_bfv_8_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_27_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_8_27_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_7_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_23_0_));
    defparam IN_MUX_bfv_7_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_24_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_7_24_0_));
    defparam IN_MUX_bfv_7_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_25_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_7_25_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_7_16_0_));
    ICE_GB \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQOU9A_0_31  (
            .USERSIGNALTOGLOBALBUFFER(N__14045),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.N_32_g ));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__12431),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_180_i_g ));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__18785),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_178_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__8372),
            .CLKHFEN(N__8374),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__8373),
            .RGB2PWM(N__8393),
            .RGB1(rgb_g),
            .CURREN(N__8387),
            .RGB2(rgb_b),
            .RGB1PWM(N__8351),
            .RGB0PWM(N__20902),
            .RGB0(rgb_r));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_0  (
            .USERSIGNALTOGLOBALBUFFER(N__15449),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_181_i_g ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__8584),
            .in2(N__8510),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__8558),
            .in2(_gnd_net_),
            .in3(N__8300),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__8531),
            .in2(N__8501),
            .in3(N__8297),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(N__9143),
            .in2(_gnd_net_),
            .in3(N__8294),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__9122),
            .in2(_gnd_net_),
            .in3(N__8291),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9098),
            .in3(N__8288),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__9074),
            .in2(_gnd_net_),
            .in3(N__8285),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9053),
            .in3(N__8282),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__9029),
            .in2(_gnd_net_),
            .in3(N__8327),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__9008),
            .in2(_gnd_net_),
            .in3(N__8324),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__8987),
            .in2(_gnd_net_),
            .in3(N__8321),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(N__9323),
            .in2(_gnd_net_),
            .in3(N__8318),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4  (
            .in0(_gnd_net_),
            .in1(N__9290),
            .in2(_gnd_net_),
            .in3(N__8315),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(N__9269),
            .in2(_gnd_net_),
            .in3(N__8312),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(N__9248),
            .in2(_gnd_net_),
            .in3(N__8309),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__9227),
            .in2(_gnd_net_),
            .in3(N__8306),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(N__9206),
            .in2(_gnd_net_),
            .in3(N__8303),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(N__9185),
            .in2(_gnd_net_),
            .in3(N__8399),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2  (
            .in0(_gnd_net_),
            .in1(N__9164),
            .in2(_gnd_net_),
            .in3(N__8396),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_0_LC_1_29_1.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_1_29_1.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_1_29_1.LUT_INIT=16'b1010101001010101;
    LogicCell40 rgb_drv_RNO_0_LC_1_29_1 (
            .in0(N__21571),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20900),
            .lcout(N_39_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_30_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_30_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_30_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_LC_1_30_2.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_1_30_2.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_1_30_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_drv_RNO_LC_1_30_2 (
            .in0(N__20901),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21575),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_16_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_16_0 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_16_0  (
            .in0(N__8649),
            .in1(N__8928),
            .in2(N__8819),
            .in3(N__8345),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21189),
            .ce(),
            .sr(N__20820));
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_2_17_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_2_17_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_2_17_1  (
            .in0(N__8927),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8621),
            .lcout(\phase_controller_slave.stoper_tr.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_1_LC_2_17_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_1_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_1_LC_2_17_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNII60D_1_LC_2_17_3  (
            .in0(N__8926),
            .in1(N__8620),
            .in2(_gnd_net_),
            .in3(N__8800),
            .lcout(\phase_controller_slave.stoper_tr.stoper_state_RNII60DZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_2_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_2_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_2_18_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_3_LC_2_18_0  (
            .in0(N__8678),
            .in1(N__8938),
            .in2(N__8336),
            .in3(N__8796),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21178),
            .ce(),
            .sr(N__20831));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_2_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_2_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_2_18_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_4_LC_2_18_1  (
            .in0(N__8793),
            .in1(N__8682),
            .in2(N__8951),
            .in3(N__8447),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21178),
            .ce(),
            .sr(N__20831));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_2_18_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_2_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_2_18_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_5_LC_2_18_2  (
            .in0(N__8679),
            .in1(N__8939),
            .in2(N__8441),
            .in3(N__8797),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21178),
            .ce(),
            .sr(N__20831));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_2_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_2_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_2_18_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_6_LC_2_18_3  (
            .in0(N__8794),
            .in1(N__8683),
            .in2(N__8952),
            .in3(N__8432),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21178),
            .ce(),
            .sr(N__20831));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_2_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_2_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_2_18_4 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_7_LC_2_18_4  (
            .in0(N__8680),
            .in1(N__8940),
            .in2(N__8426),
            .in3(N__8798),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21178),
            .ce(),
            .sr(N__20831));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_2_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_2_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_2_18_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_8_LC_2_18_5  (
            .in0(N__8795),
            .in1(N__8684),
            .in2(N__8953),
            .in3(N__8417),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21178),
            .ce(),
            .sr(N__20831));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6  (
            .in0(N__8681),
            .in1(N__8941),
            .in2(N__8411),
            .in3(N__8799),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21178),
            .ce(),
            .sr(N__20831));
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_2_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_2_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_2_19_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_0_LC_2_19_0  (
            .in0(N__9417),
            .in1(N__8669),
            .in2(N__8945),
            .in3(N__8779),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21173),
            .ce(),
            .sr(N__20837));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_2_19_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_2_19_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_2_19_1  (
            .in0(N__8773),
            .in1(N__8585),
            .in2(_gnd_net_),
            .in3(N__9416),
            .lcout(),
            .ltout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_2_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_2_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_2_19_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_1_LC_2_19_2  (
            .in0(N__8903),
            .in1(N__8668),
            .in2(N__8402),
            .in3(N__8778),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21173),
            .ce(),
            .sr(N__20837));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(N__8761),
            .in2(_gnd_net_),
            .in3(N__9414),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_2_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_2_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_2_19_4 .LUT_INIT=16'b0000010111000000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_1_LC_2_19_4  (
            .in0(N__9418),
            .in1(N__8670),
            .in2(N__8946),
            .in3(N__8780),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21173),
            .ce(),
            .sr(N__20837));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUS53_LC_2_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUS53_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUS53_LC_2_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUS53_LC_2_19_5  (
            .in0(_gnd_net_),
            .in1(N__8762),
            .in2(_gnd_net_),
            .in3(N__9415),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIUSZ0Z53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_19_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_19_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_19_6  (
            .in0(N__8902),
            .in1(N__8667),
            .in2(N__8492),
            .in3(N__8777),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21173),
            .ce(),
            .sr(N__20837));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_19_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_19_7  (
            .in0(N__8666),
            .in1(N__8904),
            .in2(N__8810),
            .in3(N__8483),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21173),
            .ce(),
            .sr(N__20837));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_20_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_20_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_20_0  (
            .in0(N__8789),
            .in1(N__8674),
            .in2(N__8947),
            .in3(N__8477),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21163),
            .ce(),
            .sr(N__20839));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_20_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_20_1 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_20_1  (
            .in0(N__8671),
            .in1(N__8911),
            .in2(N__8816),
            .in3(N__8471),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21163),
            .ce(),
            .sr(N__20839));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_20_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_20_2  (
            .in0(N__8790),
            .in1(N__8675),
            .in2(N__8948),
            .in3(N__8465),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21163),
            .ce(),
            .sr(N__20839));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_20_3 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_20_3  (
            .in0(N__8672),
            .in1(N__8912),
            .in2(N__8817),
            .in3(N__8459),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21163),
            .ce(),
            .sr(N__20839));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_20_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_20_4  (
            .in0(N__8791),
            .in1(N__8676),
            .in2(N__8949),
            .in3(N__8453),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21163),
            .ce(),
            .sr(N__20839));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_20_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_20_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_20_5  (
            .in0(N__8673),
            .in1(N__8913),
            .in2(N__8818),
            .in3(N__8966),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21163),
            .ce(),
            .sr(N__20839));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_20_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_20_6  (
            .in0(N__8792),
            .in1(N__8677),
            .in2(N__8950),
            .in3(N__8960),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21163),
            .ce(),
            .sr(N__20839));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_3_17_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_3_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_3_17_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_2_LC_3_17_0  (
            .in0(N__8648),
            .in1(N__8811),
            .in2(N__8954),
            .in3(N__8831),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21179),
            .ce(),
            .sr(N__20821));
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_3_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_3_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_3_17_4 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_LC_3_17_4  (
            .in0(N__9391),
            .in1(N__8812),
            .in2(N__8693),
            .in3(N__9422),
            .lcout(\phase_controller_slave.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21179),
            .ce(),
            .sr(N__20821));
    defparam \phase_controller_slave.start_timer_tr_LC_3_17_6 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_LC_3_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_tr_LC_3_17_6 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \phase_controller_slave.start_timer_tr_LC_3_17_6  (
            .in0(N__9362),
            .in1(N__8665),
            .in2(N__9827),
            .in3(N__9838),
            .lcout(\phase_controller_slave.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21179),
            .ce(),
            .sr(N__20821));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__9344),
            .in2(N__8567),
            .in3(N__8583),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_18_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_3_18_1  (
            .in0(N__8551),
            .in1(N__9503),
            .in2(N__8540),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_18_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_3_18_2  (
            .in0(N__8530),
            .in1(N__9350),
            .in2(N__8519),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__9329),
            .in2(N__9131),
            .in3(N__9142),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(N__9485),
            .in2(N__9107),
            .in3(N__9118),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(N__9476),
            .in2(N__9083),
            .in3(N__9094),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__9356),
            .in2(N__9062),
            .in3(N__9073),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__9338),
            .in2(N__9038),
            .in3(N__9049),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__9449),
            .in2(N__9017),
            .in3(N__9028),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__9608),
            .in2(N__8996),
            .in3(N__9007),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__9614),
            .in2(N__8975),
            .in3(N__8986),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_19_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__9599),
            .in2(N__9299),
            .in3(N__9322),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_19_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_19_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_3_19_4  (
            .in0(N__9289),
            .in1(N__9494),
            .in2(N__9278),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_19_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__9464),
            .in2(N__9257),
            .in3(N__9268),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_19_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__9455),
            .in2(N__9236),
            .in3(N__9247),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_19_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__9623),
            .in2(N__9215),
            .in3(N__9226),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_20_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__9437),
            .in2(N__9194),
            .in3(N__9205),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_20_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__9431),
            .in2(N__9173),
            .in3(N__9184),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_20_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__9593),
            .in2(N__9152),
            .in3(N__9163),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9425),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_0_LC_4_16_0 .C_ON=1'b0;
    defparam \phase_controller_slave.state_0_LC_4_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_0_LC_4_16_0 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \phase_controller_slave.state_0_LC_4_16_0  (
            .in0(N__9751),
            .in1(N__9686),
            .in2(N__9395),
            .in3(N__9374),
            .lcout(\phase_controller_slave.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21180),
            .ce(),
            .sr(N__20813));
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_4_17_0 .C_ON=1'b0;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_4_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.state_RNIVDE2_0_LC_4_17_0  (
            .in0(_gnd_net_),
            .in1(N__9390),
            .in2(_gnd_net_),
            .in3(N__9373),
            .lcout(\phase_controller_slave.state_RNIVDE2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_4_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_4_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_tr_RNO_0_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(N__9749),
            .in2(_gnd_net_),
            .in3(N__9684),
            .lcout(\phase_controller_slave.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_0 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_7_LC_4_18_0  (
            .in0(N__11874),
            .in1(N__11614),
            .in2(N__13805),
            .in3(N__11770),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21164),
            .ce(N__9575),
            .sr(N__20822));
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_3 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_3_LC_4_18_3  (
            .in0(N__11612),
            .in1(N__15113),
            .in2(N__11785),
            .in3(N__11877),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21164),
            .ce(N__9575),
            .sr(N__20822));
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_4_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_4_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_4_18_4 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_1_LC_4_18_4  (
            .in0(N__11873),
            .in1(N__11611),
            .in2(N__13544),
            .in3(N__11763),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21164),
            .ce(N__9575),
            .sr(N__20822));
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_5 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_8_LC_4_18_5  (
            .in0(N__11615),
            .in1(N__11876),
            .in2(N__11787),
            .in3(N__12630),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21164),
            .ce(N__9575),
            .sr(N__20822));
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_4_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_4_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_4_18_7 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_4_LC_4_18_7  (
            .in0(N__11613),
            .in1(N__11875),
            .in2(N__11786),
            .in3(N__15032),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21164),
            .ce(N__9575),
            .sr(N__20822));
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_4_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_4_19_0 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_4_19_0 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_2_LC_4_19_0  (
            .in0(N__14918),
            .in1(N__11202),
            .in2(N__11240),
            .in3(N__10159),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21157),
            .ce(N__9583),
            .sr(N__20827));
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_4_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_4_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_4_19_2 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_13_LC_4_19_2  (
            .in0(N__11610),
            .in1(N__11761),
            .in2(N__11900),
            .in3(N__14806),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21157),
            .ce(N__9583),
            .sr(N__20827));
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_4_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_4_19_4 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_4_19_4 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_5_LC_4_19_4  (
            .in0(N__11239),
            .in1(N__13430),
            .in2(N__11207),
            .in3(N__10160),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21157),
            .ce(N__9583),
            .sr(N__20827));
    defparam \phase_controller_slave.stoper_tr.target_timeZ0Z_6_LC_4_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_timeZ0Z_6_LC_4_19_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.stoper_tr.target_timeZ0Z_6_LC_4_19_5 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \phase_controller_slave.stoper_tr.target_timeZ0Z_6_LC_4_19_5  (
            .in0(N__13649),
            .in1(N__11893),
            .in2(N__11784),
            .in3(N__11609),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21157),
            .ce(N__9583),
            .sr(N__20827));
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_4_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_4_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_4_19_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_14_LC_4_19_7  (
            .in0(N__11762),
            .in1(N__13580),
            .in2(_gnd_net_),
            .in3(N__13727),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21157),
            .ce(N__9583),
            .sr(N__20827));
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_4_20_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_4_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_4_20_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_15_LC_4_20_0  (
            .in0(_gnd_net_),
            .in1(N__13718),
            .in2(_gnd_net_),
            .in3(N__11750),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21151),
            .ce(N__9582),
            .sr(N__20832));
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_4_20_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_4_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_4_20_1 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_9_LC_4_20_1  (
            .in0(N__11582),
            .in1(N__11781),
            .in2(N__13726),
            .in3(N__13468),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21151),
            .ce(N__9582),
            .sr(N__20832));
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_4_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_4_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_4_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_17_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13508),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21151),
            .ce(N__9582),
            .sr(N__20832));
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_4_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_4_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_4_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_18_LC_4_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15066),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21151),
            .ce(N__9582),
            .sr(N__20832));
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_4_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_4_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_4_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_16_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13760),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21151),
            .ce(N__9582),
            .sr(N__20832));
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_4_20_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_4_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_4_20_5 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_11_LC_4_20_5  (
            .in0(N__11580),
            .in1(N__14842),
            .in2(N__11782),
            .in3(N__11898),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21151),
            .ce(N__9582),
            .sr(N__20832));
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_4_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_4_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_4_20_6 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_10_LC_4_20_6  (
            .in0(N__11897),
            .in1(N__11751),
            .in2(N__14882),
            .in3(N__11579),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21151),
            .ce(N__9582),
            .sr(N__20832));
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_4_20_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_4_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_4_20_7 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_12_LC_4_20_7  (
            .in0(N__11581),
            .in1(N__13612),
            .in2(N__11783),
            .in3(N__11899),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21151),
            .ce(N__9582),
            .sr(N__20832));
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_4_21_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_4_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_4_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_19_LC_4_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16933),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21145),
            .ce(N__9587),
            .sr(N__20838));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_4_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_4_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_4_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_4_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16934),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21138),
            .ce(N__12035),
            .sr(N__20843));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_10_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_10_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_5_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9539),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21194),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_5_12_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_5_12_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_5_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_5_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9527),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21192),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_5_12_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_5_12_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_5_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_5_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9509),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21192),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_13_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_13_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_5_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9710),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21190),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_5_14_6 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_5_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_1_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__13923),
            .in2(_gnd_net_),
            .in3(N__9636),
            .lcout(\phase_controller_slave.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_5_16_1 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_5_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_0_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(N__9657),
            .in2(_gnd_net_),
            .in3(N__9864),
            .lcout(\phase_controller_slave.start_timer_hc_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_LC_5_17_0 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_LC_5_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_hc_LC_5_17_0 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \phase_controller_slave.start_timer_hc_LC_5_17_0  (
            .in0(N__9701),
            .in1(N__9692),
            .in2(N__9823),
            .in3(N__11428),
            .lcout(\phase_controller_slave.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21165),
            .ce(),
            .sr(N__20814));
    defparam \phase_controller_slave.state_1_LC_5_17_5 .C_ON=1'b0;
    defparam \phase_controller_slave.state_1_LC_5_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_1_LC_5_17_5 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_slave.state_1_LC_5_17_5  (
            .in0(N__9866),
            .in1(N__9750),
            .in2(N__9662),
            .in3(N__9685),
            .lcout(\phase_controller_slave.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21165),
            .ce(),
            .sr(N__20814));
    defparam \phase_controller_slave.state_2_LC_5_17_6 .C_ON=1'b0;
    defparam \phase_controller_slave.state_2_LC_5_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_2_LC_5_17_6 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_slave.state_2_LC_5_17_6  (
            .in0(N__9644),
            .in1(N__9658),
            .in2(N__13930),
            .in3(N__9865),
            .lcout(\phase_controller_slave.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21165),
            .ce(),
            .sr(N__20814));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_5_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_5_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_5_18_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_12_LC_5_18_5  (
            .in0(N__11427),
            .in1(N__11360),
            .in2(N__13289),
            .in3(N__10001),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21158),
            .ce(),
            .sr(N__20819));
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(N__11426),
            .in2(_gnd_net_),
            .in3(N__11359),
            .lcout(\phase_controller_slave.stoper_hc.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_3_LC_5_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.state_3_LC_5_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_3_LC_5_19_0 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \phase_controller_slave.state_3_LC_5_19_0  (
            .in0(N__9785),
            .in1(N__13916),
            .in2(N__9822),
            .in3(N__9643),
            .lcout(\phase_controller_slave.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21152),
            .ce(),
            .sr(N__20823));
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_5_19_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_5_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_5_19_1 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_LC_5_19_1  (
            .in0(N__9863),
            .in1(N__13288),
            .in2(N__9875),
            .in3(N__13145),
            .lcout(\phase_controller_slave.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21152),
            .ce(),
            .sr(N__20823));
    defparam \phase_controller_slave.state_4_LC_5_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.state_4_LC_5_19_4 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.state_4_LC_5_19_4 .LUT_INIT=16'b1100111011101110;
    LogicCell40 \phase_controller_slave.state_4_LC_5_19_4  (
            .in0(N__9812),
            .in1(N__9842),
            .in2(N__21555),
            .in3(N__9779),
            .lcout(\phase_controller_slave.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21152),
            .ce(),
            .sr(N__20823));
    defparam \phase_controller_slave.state_RNO_0_3_LC_5_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.state_RNO_0_3_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_RNO_0_3_LC_5_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.state_RNO_0_3_LC_5_20_4  (
            .in0(_gnd_net_),
            .in1(N__21556),
            .in2(_gnd_net_),
            .in3(N__9771),
            .lcout(\phase_controller_slave.state_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.T01_LC_5_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_5_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_5_21_3 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.T01_LC_5_21_3  (
            .in0(N__21487),
            .in1(N__19505),
            .in2(N__9778),
            .in3(N__15215),
            .lcout(shift_flag_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21142),
            .ce(),
            .sr(N__20833));
    defparam \phase_controller_slave.S2_LC_5_21_4 .C_ON=1'b0;
    defparam \phase_controller_slave.S2_LC_5_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S2_LC_5_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.S2_LC_5_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9755),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21142),
            .ce(),
            .sr(N__20833));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_5_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_5_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_5_24_1 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_5_24_1  (
            .in0(N__11890),
            .in1(N__14881),
            .in2(N__11788),
            .in3(N__11616),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21128),
            .ce(N__12029),
            .sr(N__20844));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_5_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_5_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_5_24_4 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_5_24_4  (
            .in0(N__11617),
            .in1(N__11777),
            .in2(N__14849),
            .in3(N__11891),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21128),
            .ce(N__12029),
            .sr(N__20844));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_5_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_5_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_5_24_7 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_5_24_7  (
            .in0(N__13725),
            .in1(N__13472),
            .in2(N__11789),
            .in3(N__11618),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21128),
            .ce(N__12029),
            .sr(N__20844));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10490),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21186),
            .ce(N__10889),
            .sr(N__20783));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10472),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21186),
            .ce(N__10889),
            .sr(N__20783));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_7_13_0  (
            .in0(N__17636),
            .in1(N__10488),
            .in2(_gnd_net_),
            .in3(N__9902),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__21181),
            .ce(N__17498),
            .sr(N__20788));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_7_13_1  (
            .in0(N__17536),
            .in1(N__10470),
            .in2(_gnd_net_),
            .in3(N__9899),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__21181),
            .ce(N__17498),
            .sr(N__20788));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_7_13_2  (
            .in0(N__17637),
            .in1(N__10449),
            .in2(_gnd_net_),
            .in3(N__9896),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__21181),
            .ce(N__17498),
            .sr(N__20788));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_7_13_3  (
            .in0(N__17537),
            .in1(N__10425),
            .in2(_gnd_net_),
            .in3(N__9893),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__21181),
            .ce(N__17498),
            .sr(N__20788));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_7_13_4  (
            .in0(N__17638),
            .in1(N__10403),
            .in2(_gnd_net_),
            .in3(N__9890),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__21181),
            .ce(N__17498),
            .sr(N__20788));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_7_13_5  (
            .in0(N__17538),
            .in1(N__10667),
            .in2(_gnd_net_),
            .in3(N__9887),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__21181),
            .ce(N__17498),
            .sr(N__20788));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_7_13_6  (
            .in0(N__17639),
            .in1(N__10647),
            .in2(_gnd_net_),
            .in3(N__9884),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__21181),
            .ce(N__17498),
            .sr(N__20788));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_7_13_7  (
            .in0(N__17539),
            .in1(N__10623),
            .in2(_gnd_net_),
            .in3(N__9881),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__21181),
            .ce(N__17498),
            .sr(N__20788));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_7_14_0  (
            .in0(N__17573),
            .in1(N__10600),
            .in2(_gnd_net_),
            .in3(N__9878),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__21174),
            .ce(N__17500),
            .sr(N__20793));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_7_14_1  (
            .in0(N__17577),
            .in1(N__10579),
            .in2(_gnd_net_),
            .in3(N__9929),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__21174),
            .ce(N__17500),
            .sr(N__20793));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_7_14_2  (
            .in0(N__17570),
            .in1(N__10557),
            .in2(_gnd_net_),
            .in3(N__9926),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__21174),
            .ce(N__17500),
            .sr(N__20793));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_7_14_3  (
            .in0(N__17574),
            .in1(N__10533),
            .in2(_gnd_net_),
            .in3(N__9923),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__21174),
            .ce(N__17500),
            .sr(N__20793));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_7_14_4  (
            .in0(N__17571),
            .in1(N__10511),
            .in2(_gnd_net_),
            .in3(N__9920),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__21174),
            .ce(N__17500),
            .sr(N__20793));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_7_14_5  (
            .in0(N__17575),
            .in1(N__10859),
            .in2(_gnd_net_),
            .in3(N__9917),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__21174),
            .ce(N__17500),
            .sr(N__20793));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_7_14_6  (
            .in0(N__17572),
            .in1(N__10839),
            .in2(_gnd_net_),
            .in3(N__9914),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__21174),
            .ce(N__17500),
            .sr(N__20793));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_7_14_7  (
            .in0(N__17576),
            .in1(N__10815),
            .in2(_gnd_net_),
            .in3(N__9911),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__21174),
            .ce(N__17500),
            .sr(N__20793));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_7_15_0  (
            .in0(N__17617),
            .in1(N__10792),
            .in2(_gnd_net_),
            .in3(N__9908),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__21166),
            .ce(N__17499),
            .sr(N__20800));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_7_15_1  (
            .in0(N__17587),
            .in1(N__10771),
            .in2(_gnd_net_),
            .in3(N__9905),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__21166),
            .ce(N__17499),
            .sr(N__20800));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_7_15_2  (
            .in0(N__17618),
            .in1(N__10749),
            .in2(_gnd_net_),
            .in3(N__9956),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__21166),
            .ce(N__17499),
            .sr(N__20800));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_7_15_3  (
            .in0(N__17588),
            .in1(N__10725),
            .in2(_gnd_net_),
            .in3(N__9953),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__21166),
            .ce(N__17499),
            .sr(N__20800));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_7_15_4  (
            .in0(N__17619),
            .in1(N__10703),
            .in2(_gnd_net_),
            .in3(N__9950),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__21166),
            .ce(N__17499),
            .sr(N__20800));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_7_15_5  (
            .in0(N__17589),
            .in1(N__10685),
            .in2(_gnd_net_),
            .in3(N__9947),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__21166),
            .ce(N__17499),
            .sr(N__20800));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_7_15_6  (
            .in0(N__17620),
            .in1(N__11052),
            .in2(_gnd_net_),
            .in3(N__9944),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__21166),
            .ce(N__17499),
            .sr(N__20800));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_7_15_7  (
            .in0(N__17590),
            .in1(N__11028),
            .in2(_gnd_net_),
            .in3(N__9941),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__21166),
            .ce(N__17499),
            .sr(N__20800));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_7_16_0  (
            .in0(N__17621),
            .in1(N__11005),
            .in2(_gnd_net_),
            .in3(N__9938),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__21159),
            .ce(N__17501),
            .sr(N__20805));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_7_16_1  (
            .in0(N__17625),
            .in1(N__10984),
            .in2(_gnd_net_),
            .in3(N__9935),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__21159),
            .ce(N__17501),
            .sr(N__20805));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_7_16_2  (
            .in0(N__17622),
            .in1(N__10950),
            .in2(_gnd_net_),
            .in3(N__9932),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__21159),
            .ce(N__17501),
            .sr(N__20805));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_7_16_3  (
            .in0(N__17626),
            .in1(N__10914),
            .in2(_gnd_net_),
            .in3(N__9980),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__21159),
            .ce(N__17501),
            .sr(N__20805));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_7_16_4  (
            .in0(N__17623),
            .in1(N__10964),
            .in2(_gnd_net_),
            .in3(N__9977),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__21159),
            .ce(N__17501),
            .sr(N__20805));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_16_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_7_16_5  (
            .in0(N__10928),
            .in1(N__17624),
            .in2(_gnd_net_),
            .in3(N__9974),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21159),
            .ce(N__17501),
            .sr(N__20805));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_17_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__13162),
            .in2(N__11063),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_7_17_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_7_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__12902),
            .in2(_gnd_net_),
            .in3(N__9971),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_7_17_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_7_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__12866),
            .in2(N__11168),
            .in3(N__9968),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_7_17_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_7_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__12833),
            .in2(_gnd_net_),
            .in3(N__9965),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_7_17_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_7_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__12803),
            .in2(_gnd_net_),
            .in3(N__9962),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_7_17_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_7_17_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12776),
            .in3(N__9959),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_7_17_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_7_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__12752),
            .in2(_gnd_net_),
            .in3(N__10016),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_7_17_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_7_17_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13085),
            .in3(N__10013),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_7_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_7_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(N__13061),
            .in2(_gnd_net_),
            .in3(N__10010),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_7_18_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_7_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_7_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(N__13040),
            .in2(_gnd_net_),
            .in3(N__10007),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_7_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_7_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(N__13019),
            .in2(_gnd_net_),
            .in3(N__10004),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_7_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_7_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(N__12998),
            .in2(_gnd_net_),
            .in3(N__9992),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_7_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_7_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(N__12971),
            .in2(_gnd_net_),
            .in3(N__9989),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_7_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_7_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(N__12950),
            .in2(_gnd_net_),
            .in3(N__9986),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_7_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_7_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(N__13397),
            .in2(_gnd_net_),
            .in3(N__9983),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_7_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_7_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(N__13376),
            .in2(_gnd_net_),
            .in3(N__10037),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_7_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_7_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__13355),
            .in2(_gnd_net_),
            .in3(N__10034),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_7_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_7_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__13334),
            .in2(_gnd_net_),
            .in3(N__10031),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_7_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_7_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__13313),
            .in2(_gnd_net_),
            .in3(N__10028),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_startlto19_LC_7_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto19_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto19_LC_7_19_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_startlto19_LC_7_19_4  (
            .in0(N__11707),
            .in1(N__11540),
            .in2(_gnd_net_),
            .in3(N__13712),
            .lcout(\phase_controller_inst1.stoper_tr.un1_start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_startlto6_LC_7_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto6_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto6_LC_7_20_0 .LUT_INIT=16'b1010100010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_startlto6_LC_7_20_0  (
            .in0(N__13641),
            .in1(N__14906),
            .in2(N__15112),
            .in3(N__10022),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un1_startlt8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_startlto9_0_0_LC_7_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto9_0_0_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto9_0_0_LC_7_20_1 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_startlto9_0_0_LC_7_20_1  (
            .in0(N__13575),
            .in1(N__13467),
            .in2(N__10025),
            .in3(N__11249),
            .lcout(\phase_controller_inst1.stoper_tr.un1_startlt15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_startlto5_1_LC_7_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto5_1_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto5_1_LC_7_20_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_startlto5_1_LC_7_20_3  (
            .in0(N__13418),
            .in1(N__13530),
            .in2(_gnd_net_),
            .in3(N__15020),
            .lcout(\phase_controller_inst1.stoper_tr.un1_startlto5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_4_LC_7_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_4_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_4_LC_7_20_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un2_startlto19_4_LC_7_20_4  (
            .in0(N__15056),
            .in1(N__16925),
            .in2(_gnd_net_),
            .in3(N__13691),
            .lcout(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un2_startlto6_0_LC_7_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto6_0_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto6_0_LC_7_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un2_startlto6_0_LC_7_20_5  (
            .in0(N__13419),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13640),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un2_startlto6Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un2_startlto6_LC_7_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto6_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto6_LC_7_20_6 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un2_startlto6_LC_7_20_6  (
            .in0(N__15021),
            .in1(N__15107),
            .in2(N__10049),
            .in3(N__14907),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un2_startlt19_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_9_LC_7_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_9_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_9_LC_7_20_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un2_startlto19_9_LC_7_20_7  (
            .in0(N__10046),
            .in1(N__13611),
            .in2(N__10040),
            .in3(N__14841),
            .lcout(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_7_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_7_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_7_21_2 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_7_21_2  (
            .in0(N__11838),
            .in1(N__11541),
            .in2(N__14807),
            .in3(N__11675),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21133),
            .ce(N__12031),
            .sr(N__20824));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_7_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_7_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_7_21_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(N__11674),
            .in2(_gnd_net_),
            .in3(N__13713),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21133),
            .ce(N__12031),
            .sr(N__20824));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_22_0 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_22_0 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_7_22_0  (
            .in0(N__10158),
            .in1(N__11226),
            .in2(N__11206),
            .in3(N__13426),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21129),
            .ce(N__12030),
            .sr(N__20828));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_7_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_7_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_7_22_1 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_7_22_1  (
            .in0(N__11576),
            .in1(N__11701),
            .in2(N__11872),
            .in3(N__13613),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21129),
            .ce(N__12030),
            .sr(N__20828));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_7_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_7_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_7_22_2 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_7_22_2  (
            .in0(N__15111),
            .in1(N__11843),
            .in2(N__11749),
            .in3(N__11578),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21129),
            .ce(N__12030),
            .sr(N__20828));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_7_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_7_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_7_22_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_7_22_3  (
            .in0(N__11706),
            .in1(N__13579),
            .in2(_gnd_net_),
            .in3(N__13714),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21129),
            .ce(N__12030),
            .sr(N__20828));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_7_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_7_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_7_22_4 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_7_22_4  (
            .in0(N__11702),
            .in1(N__13537),
            .in2(N__11892),
            .in3(N__11577),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21129),
            .ce(N__12030),
            .sr(N__20828));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_7_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_7_22_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_7_22_5 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_7_22_5  (
            .in0(N__14914),
            .in1(N__11198),
            .in2(N__11230),
            .in3(N__10157),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21129),
            .ce(N__12030),
            .sr(N__20828));
    defparam \phase_controller_inst1.stoper_tr.target_timeZ0Z_6_LC_7_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_timeZ0Z_6_LC_7_22_6 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.stoper_tr.target_timeZ0Z_6_LC_7_22_6 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_timeZ0Z_6_LC_7_22_6  (
            .in0(N__13648),
            .in1(N__11842),
            .in2(N__11748),
            .in3(N__11575),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21129),
            .ce(N__12030),
            .sr(N__20828));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_7_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_7_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_7_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_7_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15071),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21129),
            .ce(N__12030),
            .sr(N__20828));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__10136),
            .in2(N__10130),
            .in3(N__11973),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_7_23_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_23_1  (
            .in0(_gnd_net_),
            .in1(N__10121),
            .in2(N__10115),
            .in3(N__11947),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_23_2  (
            .in0(_gnd_net_),
            .in1(N__10106),
            .in2(N__10100),
            .in3(N__12205),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_23_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_23_3  (
            .in0(_gnd_net_),
            .in1(N__11936),
            .in2(N__10091),
            .in3(N__12169),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_23_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_23_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(N__10082),
            .in2(N__10076),
            .in3(N__12148),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_23_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_23_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_23_5  (
            .in0(_gnd_net_),
            .in1(N__10067),
            .in2(N__10058),
            .in3(N__12127),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_23_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_23_6  (
            .in0(_gnd_net_),
            .in1(N__11507),
            .in2(N__10295),
            .in3(N__12106),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_23_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_23_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_23_7  (
            .in0(_gnd_net_),
            .in1(N__11918),
            .in2(N__10286),
            .in3(N__12082),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_24_0  (
            .in0(_gnd_net_),
            .in1(N__10277),
            .in2(N__10268),
            .in3(N__12058),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_7_24_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_24_1  (
            .in0(_gnd_net_),
            .in1(N__10259),
            .in2(N__10247),
            .in3(N__12397),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_24_2  (
            .in0(_gnd_net_),
            .in1(N__10238),
            .in2(N__10229),
            .in3(N__12371),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_24_3  (
            .in0(_gnd_net_),
            .in1(N__10220),
            .in2(N__10208),
            .in3(N__13955),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_24_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_24_4  (
            .in0(_gnd_net_),
            .in1(N__10199),
            .in2(N__10190),
            .in3(N__12344),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_24_5  (
            .in0(_gnd_net_),
            .in1(N__10181),
            .in2(N__10169),
            .in3(N__12319),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_24_6  (
            .in0(_gnd_net_),
            .in1(N__10376),
            .in2(N__10364),
            .in3(N__12290),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_24_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_24_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_24_7  (
            .in0(_gnd_net_),
            .in1(N__11912),
            .in2(N__10355),
            .in3(N__12266),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_25_0  (
            .in0(_gnd_net_),
            .in1(N__11930),
            .in2(N__10346),
            .in3(N__12238),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_7_25_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_25_1  (
            .in0(_gnd_net_),
            .in1(N__10337),
            .in2(N__10328),
            .in3(N__12472),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_25_2  (
            .in0(_gnd_net_),
            .in1(N__10319),
            .in2(N__10307),
            .in3(N__12451),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10298),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_7_25_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_7_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_7_25_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_7_25_4  (
            .in0(N__15853),
            .in1(_gnd_net_),
            .in2(N__15935),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_25_5  (
            .in0(_gnd_net_),
            .in1(N__15852),
            .in2(_gnd_net_),
            .in3(N__15922),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_25_6 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_25_6  (
            .in0(N__15854),
            .in1(_gnd_net_),
            .in2(N__11984),
            .in3(N__15926),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_26_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_26_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_26_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_26_0  (
            .in0(N__15883),
            .in1(N__15587),
            .in2(N__15740),
            .in3(N__12329),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(N__20845));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_26_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_26_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_26_1 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_26_1  (
            .in0(N__15588),
            .in1(N__15729),
            .in2(N__12302),
            .in3(N__15887),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(N__20845));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_26_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_26_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_26_2  (
            .in0(N__15884),
            .in1(N__15589),
            .in2(N__15741),
            .in3(N__12275),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(N__20845));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_26_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_26_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_26_3 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_26_3  (
            .in0(N__15590),
            .in1(N__15730),
            .in2(N__12251),
            .in3(N__15888),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(N__20845));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_26_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_26_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_26_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_26_4  (
            .in0(N__15885),
            .in1(N__15591),
            .in2(N__15742),
            .in3(N__12227),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(N__20845));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_26_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_26_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_26_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_26_5  (
            .in0(N__15592),
            .in1(N__15731),
            .in2(N__15899),
            .in3(N__12461),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(N__20845));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_26_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_26_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_26_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_26_6  (
            .in0(N__15886),
            .in1(N__15593),
            .in2(N__15743),
            .in3(N__12437),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(N__20845));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_26_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_26_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_26_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_26_7  (
            .in0(N__15586),
            .in1(N__15728),
            .in2(N__15898),
            .in3(N__12356),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(N__20845));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_9_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_9_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10385),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21193),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_12_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_12_1  (
            .in0(N__14005),
            .in1(N__14056),
            .in2(_gnd_net_),
            .in3(N__14341),
            .lcout(\delay_measurement_inst.N_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_12_2  (
            .in0(N__17854),
            .in1(N__17734),
            .in2(N__14326),
            .in3(N__13972),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_105 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_9_LC_8_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_9_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_9_LC_8_12_3 .LUT_INIT=16'b0001000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4TEU1_9_LC_8_12_3  (
            .in0(N__18031),
            .in1(N__14082),
            .in2(N__10493),
            .in3(N__14116),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_4_LC_8_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_4_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_4_LC_8_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_4_LC_8_12_5  (
            .in0(N__12667),
            .in1(N__14182),
            .in2(N__12698),
            .in3(N__14410),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__10489),
            .in2(N__10450),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__21175),
            .ce(N__10888),
            .sr(N__20784));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__10471),
            .in2(N__10426),
            .in3(N__10454),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__21175),
            .ce(N__10888),
            .sr(N__20784));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__10401),
            .in2(N__10451),
            .in3(N__10430),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__21175),
            .ce(N__10888),
            .sr(N__20784));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__10665),
            .in2(N__10427),
            .in3(N__10406),
            .lcout(\delay_measurement_inst.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__21175),
            .ce(N__10888),
            .sr(N__20784));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__10402),
            .in2(N__10648),
            .in3(N__10388),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__21175),
            .ce(N__10888),
            .sr(N__20784));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__10666),
            .in2(N__10624),
            .in3(N__10652),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__21175),
            .ce(N__10888),
            .sr(N__20784));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__10599),
            .in2(N__10649),
            .in3(N__10628),
            .lcout(\delay_measurement_inst.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__21175),
            .ce(N__10888),
            .sr(N__20784));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__10578),
            .in2(N__10625),
            .in3(N__10604),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__21175),
            .ce(N__10888),
            .sr(N__20784));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__10601),
            .in2(N__10558),
            .in3(N__10583),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__21167),
            .ce(N__10887),
            .sr(N__20789));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__10580),
            .in2(N__10534),
            .in3(N__10562),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__21167),
            .ce(N__10887),
            .sr(N__20789));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__10509),
            .in2(N__10559),
            .in3(N__10538),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__21167),
            .ce(N__10887),
            .sr(N__20789));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__10857),
            .in2(N__10535),
            .in3(N__10514),
            .lcout(\delay_measurement_inst.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__21167),
            .ce(N__10887),
            .sr(N__20789));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__10510),
            .in2(N__10840),
            .in3(N__10496),
            .lcout(\delay_measurement_inst.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__21167),
            .ce(N__10887),
            .sr(N__20789));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__10858),
            .in2(N__10816),
            .in3(N__10844),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__21167),
            .ce(N__10887),
            .sr(N__20789));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__10791),
            .in2(N__10841),
            .in3(N__10820),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__21167),
            .ce(N__10887),
            .sr(N__20789));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__10770),
            .in2(N__10817),
            .in3(N__10796),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__21167),
            .ce(N__10887),
            .sr(N__20789));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__10793),
            .in2(N__10750),
            .in3(N__10775),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__21160),
            .ce(N__10886),
            .sr(N__20794));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__10772),
            .in2(N__10726),
            .in3(N__10754),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__21160),
            .ce(N__10886),
            .sr(N__20794));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__10701),
            .in2(N__10751),
            .in3(N__10730),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__21160),
            .ce(N__10886),
            .sr(N__20794));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__10683),
            .in2(N__10727),
            .in3(N__10706),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__21160),
            .ce(N__10886),
            .sr(N__20794));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__10702),
            .in2(N__11053),
            .in3(N__10688),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__21160),
            .ce(N__10886),
            .sr(N__20794));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__10684),
            .in2(N__11029),
            .in3(N__10670),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__21160),
            .ce(N__10886),
            .sr(N__20794));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__11004),
            .in2(N__11054),
            .in3(N__11033),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__21160),
            .ce(N__10886),
            .sr(N__20794));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__10983),
            .in2(N__11030),
            .in3(N__11009),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__21160),
            .ce(N__10886),
            .sr(N__20794));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__11006),
            .in2(N__10951),
            .in3(N__10988),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__21153),
            .ce(N__10885),
            .sr(N__20801));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(N__10985),
            .in2(N__10915),
            .in3(N__10967),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__21153),
            .ce(N__10885),
            .sr(N__20801));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(N__10963),
            .in2(N__10952),
            .in3(N__10931),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__21153),
            .ce(N__10885),
            .sr(N__20801));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(N__10927),
            .in2(N__10916),
            .in3(N__10895),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__21153),
            .ce(N__10885),
            .sr(N__20801));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10892),
            .lcout(\delay_measurement_inst.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21153),
            .ce(N__10885),
            .sr(N__20801));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_8_17_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_8_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_8_17_0 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_3_LC_8_17_0  (
            .in0(N__13281),
            .in1(N__11461),
            .in2(N__10868),
            .in3(N__11322),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(),
            .sr(N__20806));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_8_17_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_8_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_8_17_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_4_LC_8_17_1  (
            .in0(N__11458),
            .in1(N__13285),
            .in2(N__11356),
            .in3(N__11108),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(),
            .sr(N__20806));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_8_17_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_8_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_8_17_2 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_5_LC_8_17_2  (
            .in0(N__13282),
            .in1(N__11462),
            .in2(N__11102),
            .in3(N__11323),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(),
            .sr(N__20806));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_8_17_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_8_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_8_17_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_6_LC_8_17_3  (
            .in0(N__11459),
            .in1(N__13286),
            .in2(N__11357),
            .in3(N__11093),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(),
            .sr(N__20806));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_8_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_8_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_8_17_4 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_7_LC_8_17_4  (
            .in0(N__13283),
            .in1(N__11463),
            .in2(N__11087),
            .in3(N__11324),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(),
            .sr(N__20806));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_8_17_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_8_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_8_17_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_8_LC_8_17_5  (
            .in0(N__11460),
            .in1(N__13287),
            .in2(N__11358),
            .in3(N__11078),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(),
            .sr(N__20806));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_8_17_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_8_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_8_17_6 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_9_LC_8_17_6  (
            .in0(N__13284),
            .in1(N__11464),
            .in2(N__11072),
            .in3(N__11325),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(),
            .sr(N__20806));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_1_LC_8_17_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_1_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_1_LC_8_17_7 .LUT_INIT=16'b0000010000000100;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_1_LC_8_17_7  (
            .in0(N__11312),
            .in1(N__11429),
            .in2(N__13274),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.stoper_state_RNI10KLZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_8_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_8_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_8_18_0 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_1_LC_8_18_0  (
            .in0(N__13228),
            .in1(N__11466),
            .in2(N__13115),
            .in3(N__11337),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20809));
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_8_18_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_8_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_8_18_2 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_0_LC_8_18_2  (
            .in0(N__13139),
            .in1(N__11332),
            .in2(N__13271),
            .in3(N__11468),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20809));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__13225),
            .in2(_gnd_net_),
            .in3(N__13137),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_8_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_8_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_8_18_4 .LUT_INIT=16'b0001110000010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_1_LC_8_18_4  (
            .in0(N__13140),
            .in1(N__11333),
            .in2(N__13272),
            .in3(N__11469),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20809));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DK_LC_8_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DK_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DK_LC_8_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DK_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__13226),
            .in2(_gnd_net_),
            .in3(N__13138),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNI89DKZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_8_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_8_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_8_18_6 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_10_LC_8_18_6  (
            .in0(N__13227),
            .in1(N__11331),
            .in2(N__11159),
            .in3(N__11467),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20809));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_8_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_8_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_8_18_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_11_LC_8_18_7  (
            .in0(N__11465),
            .in1(N__13229),
            .in2(N__11361),
            .in3(N__11150),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20809));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_8_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_8_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_8_19_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_13_LC_8_19_0  (
            .in0(N__13248),
            .in1(N__11474),
            .in2(N__11362),
            .in3(N__11144),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21139),
            .ce(),
            .sr(N__20810));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_8_19_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_8_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_8_19_1 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_14_LC_8_19_1  (
            .in0(N__11470),
            .in1(N__13252),
            .in2(N__11138),
            .in3(N__11350),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21139),
            .ce(),
            .sr(N__20810));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_8_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_8_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_8_19_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_15_LC_8_19_2  (
            .in0(N__13249),
            .in1(N__11475),
            .in2(N__11363),
            .in3(N__11129),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21139),
            .ce(),
            .sr(N__20810));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_8_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_8_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_8_19_3 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_16_LC_8_19_3  (
            .in0(N__11471),
            .in1(N__13253),
            .in2(N__11123),
            .in3(N__11351),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21139),
            .ce(),
            .sr(N__20810));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_8_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_8_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_8_19_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_17_LC_8_19_4  (
            .in0(N__13250),
            .in1(N__11476),
            .in2(N__11364),
            .in3(N__11114),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21139),
            .ce(),
            .sr(N__20810));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_8_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_8_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_8_19_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_18_LC_8_19_5  (
            .in0(N__11472),
            .in1(N__13254),
            .in2(N__11366),
            .in3(N__11489),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21139),
            .ce(),
            .sr(N__20810));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_8_19_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_8_19_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_19_LC_8_19_6  (
            .in0(N__13251),
            .in1(N__11477),
            .in2(N__11365),
            .in3(N__11483),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21139),
            .ce(),
            .sr(N__20810));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_8_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_8_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_8_19_7 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_2_LC_8_19_7  (
            .in0(N__11473),
            .in1(N__13255),
            .in2(N__11378),
            .in3(N__11352),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21139),
            .ce(),
            .sr(N__20810));
    defparam \phase_controller_inst1.stoper_tr.un1_startlto9_c_LC_8_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto9_c_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto9_c_LC_8_20_3 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_startlto9_c_LC_8_20_3  (
            .in0(N__13456),
            .in1(N__12623),
            .in2(_gnd_net_),
            .in3(N__13794),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un1_startlto9_cZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_startlto13_3_LC_8_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto13_3_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto13_3_LC_8_20_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_startlto13_3_LC_8_20_4  (
            .in0(N__13601),
            .in1(N__14837),
            .in2(N__11252),
            .in3(N__13816),
            .lcout(\phase_controller_inst1.stoper_tr.un1_startlto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_6_LC_8_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_6_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_6_LC_8_21_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un2_startlto19_6_LC_8_21_4  (
            .in0(N__12631),
            .in1(N__13457),
            .in2(N__13798),
            .in3(N__13557),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_8_LC_8_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_8_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_8_LC_8_21_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un2_startlto19_8_LC_8_21_5  (
            .in0(N__13753),
            .in1(N__13496),
            .in2(N__11243),
            .in3(N__13817),
            .lcout(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8 ),
            .ltout(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_start_0_LC_8_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_start_0_LC_8_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_start_0_LC_8_21_6 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_start_0_LC_8_21_6  (
            .in0(N__11673),
            .in1(N__13687),
            .in2(N__11210),
            .in3(N__11181),
            .lcout(\phase_controller_inst1.stoper_tr.un3_start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_startlto19_2_LC_8_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto19_2_LC_8_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_startlto19_2_LC_8_21_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_startlto19_2_LC_8_21_7  (
            .in0(N__13752),
            .in1(N__16926),
            .in2(N__13503),
            .in3(N__15067),
            .lcout(\phase_controller_inst1.stoper_tr.un1_startlto19Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_8_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_8_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_8_22_0 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_8_22_0  (
            .in0(N__11839),
            .in1(N__15028),
            .in2(N__11745),
            .in3(N__11583),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21125),
            .ce(N__12016),
            .sr(N__20825));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_8_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_8_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_8_22_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_8_22_3  (
            .in0(N__13504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21125),
            .ce(N__12016),
            .sr(N__20825));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_8_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_8_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_8_22_4 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_8_22_4  (
            .in0(N__11841),
            .in1(N__12632),
            .in2(N__11747),
            .in3(N__11585),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21125),
            .ce(N__12016),
            .sr(N__20825));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_8_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_8_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_8_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_8_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13748),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21125),
            .ce(N__12016),
            .sr(N__20825));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_8_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_8_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_8_22_6 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_8_22_6  (
            .in0(N__11840),
            .in1(N__13792),
            .in2(N__11746),
            .in3(N__11584),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21125),
            .ce(N__12016),
            .sr(N__20825));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_23_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_23_0  (
            .in0(N__15560),
            .in1(N__15713),
            .in2(N__11501),
            .in3(N__15851),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21119),
            .ce(),
            .sr(N__20829));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_23_2 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_23_2  (
            .in0(N__15562),
            .in1(N__15714),
            .in2(N__15897),
            .in3(N__15936),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21119),
            .ce(),
            .sr(N__20829));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_23_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_23_6  (
            .in0(N__15559),
            .in1(N__15712),
            .in2(N__12386),
            .in3(N__15850),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21119),
            .ce(),
            .sr(N__20829));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_23_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_23_7  (
            .in0(N__15849),
            .in1(N__15561),
            .in2(N__15739),
            .in3(N__12218),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21119),
            .ce(),
            .sr(N__20829));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_24_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_24_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_24_0  (
            .in0(N__15828),
            .in1(N__15552),
            .in2(N__15735),
            .in3(N__12179),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21114),
            .ce(),
            .sr(N__20834));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_24_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_24_1  (
            .in0(N__15553),
            .in1(N__15832),
            .in2(N__15732),
            .in3(N__12158),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21114),
            .ce(),
            .sr(N__20834));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_24_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_24_2  (
            .in0(N__15829),
            .in1(N__15554),
            .in2(N__15736),
            .in3(N__12137),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21114),
            .ce(),
            .sr(N__20834));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_24_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_24_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_24_3  (
            .in0(N__15555),
            .in1(N__15833),
            .in2(N__15733),
            .in3(N__12116),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21114),
            .ce(),
            .sr(N__20834));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_24_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_24_4  (
            .in0(N__15830),
            .in1(N__15556),
            .in2(N__15737),
            .in3(N__12095),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21114),
            .ce(),
            .sr(N__20834));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_24_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_24_5  (
            .in0(N__15557),
            .in1(N__15834),
            .in2(N__15734),
            .in3(N__12071),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21114),
            .ce(),
            .sr(N__20834));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_24_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_24_6  (
            .in0(N__15831),
            .in1(N__15558),
            .in2(N__15738),
            .in3(N__12047),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21114),
            .ce(),
            .sr(N__20834));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_1_LC_8_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_1_LC_8_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_1_LC_8_24_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_1_LC_8_24_7  (
            .in0(N__15687),
            .in1(N__15550),
            .in2(_gnd_net_),
            .in3(N__15827),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_RNIEUJMZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_25_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_25_0  (
            .in0(_gnd_net_),
            .in1(N__11980),
            .in2(N__11960),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_25_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_25_1  (
            .in0(_gnd_net_),
            .in1(N__11951),
            .in2(_gnd_net_),
            .in3(N__12209),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_25_2  (
            .in0(_gnd_net_),
            .in1(N__12206),
            .in2(N__12188),
            .in3(N__12173),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_25_3  (
            .in0(_gnd_net_),
            .in1(N__12170),
            .in2(_gnd_net_),
            .in3(N__12152),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_25_4  (
            .in0(_gnd_net_),
            .in1(N__12149),
            .in2(_gnd_net_),
            .in3(N__12131),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_25_5  (
            .in0(_gnd_net_),
            .in1(N__12128),
            .in2(_gnd_net_),
            .in3(N__12110),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_25_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_25_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_25_6  (
            .in0(_gnd_net_),
            .in1(N__12107),
            .in2(_gnd_net_),
            .in3(N__12089),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_25_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_25_7  (
            .in0(_gnd_net_),
            .in1(N__12086),
            .in2(_gnd_net_),
            .in3(N__12065),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_26_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_26_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_26_0  (
            .in0(_gnd_net_),
            .in1(N__12062),
            .in2(_gnd_net_),
            .in3(N__12038),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_8_26_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_26_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_26_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_26_1  (
            .in0(_gnd_net_),
            .in1(N__12401),
            .in2(_gnd_net_),
            .in3(N__12374),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_26_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_26_2  (
            .in0(_gnd_net_),
            .in1(N__12370),
            .in2(_gnd_net_),
            .in3(N__12350),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_26_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_26_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_26_3  (
            .in0(_gnd_net_),
            .in1(N__13951),
            .in2(_gnd_net_),
            .in3(N__12347),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_26_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_26_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_26_4  (
            .in0(_gnd_net_),
            .in1(N__12343),
            .in2(_gnd_net_),
            .in3(N__12323),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_26_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_26_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_26_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12320),
            .in3(N__12293),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_26_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_26_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_26_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_26_6  (
            .in0(_gnd_net_),
            .in1(N__12289),
            .in2(_gnd_net_),
            .in3(N__12269),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_26_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_26_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_26_7  (
            .in0(_gnd_net_),
            .in1(N__12265),
            .in2(_gnd_net_),
            .in3(N__12242),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_27_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_27_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_27_0  (
            .in0(_gnd_net_),
            .in1(N__12239),
            .in2(_gnd_net_),
            .in3(N__12221),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_8_27_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_27_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_27_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_27_1  (
            .in0(_gnd_net_),
            .in1(N__12473),
            .in2(_gnd_net_),
            .in3(N__12455),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_27_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_27_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_27_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_27_2  (
            .in0(_gnd_net_),
            .in1(N__12452),
            .in2(_gnd_net_),
            .in3(N__12440),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_9_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_9_9_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_9_9_2  (
            .in0(N__20892),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13850),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21191),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__15477),
            .in2(_gnd_net_),
            .in3(N__17039),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_180_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_9_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_9_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_9_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_9_9_7 (
            .in0(N__12410),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21191),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_sync_1_LC_9_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_sync_1_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_sync_1_LC_9_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.tr_sync_1_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18857),
            .lcout(\delay_measurement_inst.tr_syncZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21187),
            .ce(),
            .sr(N__20769));
    defparam \delay_measurement_inst.tr_prev_LC_9_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_prev_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_prev_LC_9_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.tr_prev_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13883),
            .lcout(\delay_measurement_inst.tr_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21187),
            .ce(),
            .sr(N__20769));
    defparam \delay_measurement_inst.tr_state_0_LC_9_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_9_11_0 .LUT_INIT=16'b0000110000000110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_9_11_0  (
            .in0(N__13881),
            .in1(N__14167),
            .in2(N__20903),
            .in3(N__14152),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21182),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_RNIVV8G_0_LC_9_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_RNIVV8G_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.tr_state_RNIVV8G_0_LC_9_11_4 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \delay_measurement_inst.tr_state_RNIVV8G_0_LC_9_11_4  (
            .in0(N__13880),
            .in1(N__14166),
            .in2(_gnd_net_),
            .in3(N__14151),
            .lcout(\delay_measurement_inst.tr_state_RNIVV8GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJQC01_31_LC_9_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJQC01_31_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJQC01_31_LC_9_11_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJQC01_31_LC_9_11_6  (
            .in0(N__20894),
            .in1(N__17794),
            .in2(_gnd_net_),
            .in3(N__15381),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_9_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_9_12_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_9_12_0  (
            .in0(N__14365),
            .in1(N__12696),
            .in2(N__12671),
            .in3(N__14397),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_81 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_9_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_9_12_1 .LUT_INIT=16'b1010101011111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE5L06_31_LC_9_12_1  (
            .in0(N__17798),
            .in1(N__12533),
            .in2(N__12527),
            .in3(N__17962),
            .lcout(\delay_measurement_inst.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_9_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_9_12_2 .LUT_INIT=16'b1011101110111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBM7A4_14_LC_9_12_2  (
            .in0(N__17961),
            .in1(N__15400),
            .in2(N__18039),
            .in3(N__14115),
            .lcout(\delay_measurement_inst.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40E01_17_LC_9_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40E01_17_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40E01_17_LC_9_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40E01_17_LC_9_12_3  (
            .in0(N__14114),
            .in1(N__14364),
            .in2(N__14399),
            .in3(N__18024),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKF324_15_LC_9_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKF324_15_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKF324_15_LC_9_12_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKF324_15_LC_9_12_4  (
            .in0(N__17963),
            .in1(_gnd_net_),
            .in2(N__18038),
            .in3(N__12509),
            .lcout(\delay_measurement_inst.N_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE9BL2_2_LC_9_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE9BL2_2_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE9BL2_2_LC_9_12_5 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE9BL2_2_LC_9_12_5  (
            .in0(N__12643),
            .in1(N__12487),
            .in2(N__14086),
            .in3(N__12524),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJTHF5_17_LC_9_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJTHF5_17_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJTHF5_17_LC_9_12_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJTHF5_17_LC_9_12_6  (
            .in0(N__15388),
            .in1(N__14279),
            .in2(N__12518),
            .in3(N__12515),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_reset_1_i_a2_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQOU9A_31_LC_9_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQOU9A_31_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQOU9A_31_LC_9_12_7 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQOU9A_31_LC_9_12_7  (
            .in0(N__12508),
            .in1(N__12500),
            .in2(N__12494),
            .in3(N__17960),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_esr_2_LC_9_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_2_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_2_LC_9_13_0 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_2_LC_9_13_0  (
            .in0(N__14283),
            .in1(N__14253),
            .in2(N__14223),
            .in3(N__12491),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21168),
            .ce(N__17686),
            .sr(N__17658));
    defparam \delay_measurement_inst.delay_hc_reg_esr_19_LC_9_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_19_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_19_LC_9_13_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_19_LC_9_13_2  (
            .in0(N__17965),
            .in1(N__17796),
            .in2(_gnd_net_),
            .in3(N__12697),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21168),
            .ce(N__17686),
            .sr(N__17658));
    defparam \delay_measurement_inst.delay_hc_reg_esr_16_LC_9_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_16_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_16_LC_9_13_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_16_LC_9_13_3  (
            .in0(N__17795),
            .in1(N__17964),
            .in2(_gnd_net_),
            .in3(N__12666),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21168),
            .ce(N__17686),
            .sr(N__17658));
    defparam \delay_measurement_inst.delay_hc_reg_ess_3_LC_9_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_ess_3_LC_9_13_7 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_ess_3_LC_9_13_7 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_ess_3_LC_9_13_7  (
            .in0(N__14254),
            .in1(N__12644),
            .in2(N__14303),
            .in3(N__14211),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21168),
            .ce(N__17686),
            .sr(N__17658));
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_9_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_9_14_1 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_8_LC_9_14_1  (
            .in0(N__14996),
            .in1(N__19850),
            .in2(N__15332),
            .in3(N__12611),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21161),
            .ce(),
            .sr(N__17185));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_5  (
            .in0(N__12587),
            .in1(N__12581),
            .in2(N__12575),
            .in3(N__12566),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_7_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16261),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21154),
            .ce(N__18772),
            .sr(N__20790));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16195),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21154),
            .ce(N__18772),
            .sr(N__20790));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16166),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21154),
            .ce(N__18772),
            .sr(N__20790));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_9_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_9_15_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_9_15_4  (
            .in0(N__12560),
            .in1(N__12554),
            .in2(N__12548),
            .in3(N__12539),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_9_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_9_15_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_9_15_5  (
            .in0(N__12731),
            .in1(N__12725),
            .in2(N__12719),
            .in3(N__12704),
            .lcout(\delay_measurement_inst.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_9_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_9_15_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI23AG_29_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__12716),
            .in2(_gnd_net_),
            .in3(N__12710),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_5_0_o2_0_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16228),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21154),
            .ce(N__18772),
            .sr(N__20790));
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_9_16_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_9_16_0 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_9_16_0 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_9_16_0  (
            .in0(N__16846),
            .in1(N__16609),
            .in2(N__16442),
            .in3(N__16717),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__15141),
            .sr(N__20795));
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_9_16_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_9_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_9_16_1 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_4_LC_9_16_1  (
            .in0(N__16720),
            .in1(N__16436),
            .in2(N__16622),
            .in3(N__17362),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__15141),
            .sr(N__20795));
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_9_16_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_9_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_9_16_2 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_8_LC_9_16_2  (
            .in0(N__16437),
            .in1(N__16610),
            .in2(N__16106),
            .in3(N__16721),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__15141),
            .sr(N__20795));
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_9_16_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_9_16_3 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_9_16_3 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_2_LC_9_16_3  (
            .in0(N__17453),
            .in1(N__17238),
            .in2(N__16016),
            .in3(N__16132),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__15141),
            .sr(N__20795));
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_9_16_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_9_16_4 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_9_16_4 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_5_LC_9_16_4  (
            .in0(N__16133),
            .in1(N__16015),
            .in2(N__17243),
            .in3(N__16289),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__15141),
            .sr(N__20795));
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_9_16_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_9_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_9_16_5 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_1_LC_9_16_5  (
            .in0(N__16718),
            .in1(N__16434),
            .in2(N__16620),
            .in3(N__15980),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__15141),
            .sr(N__20795));
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_9_16_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_9_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_9_16_7 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_3_LC_9_16_7  (
            .in0(N__16719),
            .in1(N__16435),
            .in2(N__16621),
            .in3(N__17399),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__15141),
            .sr(N__20795));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_17_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__12929),
            .in2(N__12920),
            .in3(N__13161),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_17_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__12911),
            .in2(N__12884),
            .in3(N__12901),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_17_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__12875),
            .in2(N__12851),
            .in3(N__12862),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_17_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__12842),
            .in2(N__12821),
            .in3(N__12832),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_17_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__12812),
            .in2(N__12791),
            .in3(N__12802),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_17_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__12782),
            .in2(N__12761),
            .in3(N__12772),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_17_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__14756),
            .in2(N__12740),
            .in3(N__12751),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_17_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__13094),
            .in2(N__13070),
            .in3(N__13081),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__14750),
            .in2(N__13049),
            .in3(N__13060),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__14744),
            .in2(N__13028),
            .in3(N__13039),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__14765),
            .in2(N__13007),
            .in3(N__13018),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__14609),
            .in2(N__12980),
            .in3(N__12997),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__15149),
            .in2(N__12959),
            .in3(N__12970),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__14726),
            .in2(N__12938),
            .in3(N__12949),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__14735),
            .in2(N__13385),
            .in3(N__13396),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__14717),
            .in2(N__13364),
            .in3(N__13375),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__14708),
            .in2(N__13343),
            .in3(N__13354),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__14702),
            .in2(N__13322),
            .in3(N__13333),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__14603),
            .in2(N__13301),
            .in3(N__13312),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13292),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_9_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_9_19_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_9_19_5  (
            .in0(N__13273),
            .in1(N__13163),
            .in2(_gnd_net_),
            .in3(N__13141),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_9_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_9_19_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_9_19_6  (
            .in0(N__19021),
            .in1(N__19843),
            .in2(_gnd_net_),
            .in3(N__19891),
            .lcout(\delay_measurement_inst.N_172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_9_19_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_9_19_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_9_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_9_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13106),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21134),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_20_0 .LUT_INIT=16'b0000000011010000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_15_LC_9_20_0  (
            .in0(N__16980),
            .in1(N__21679),
            .in2(N__20261),
            .in3(N__15343),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(N__16892),
            .sr(N__17179));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_20_1 .LUT_INIT=16'b0010001110101111;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_9_20_1  (
            .in0(N__19025),
            .in1(N__15280),
            .in2(N__14995),
            .in3(N__14946),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(N__16892),
            .sr(N__17179));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_20_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_20_2 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_9_20_2  (
            .in0(N__21670),
            .in1(N__19657),
            .in2(_gnd_net_),
            .in3(N__15364),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(N__16892),
            .sr(N__17179));
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_20_3 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_14_LC_9_20_3  (
            .in0(N__19556),
            .in1(N__21671),
            .in2(N__15344),
            .in3(N__16982),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(N__16892),
            .sr(N__17179));
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_20_4 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_20_4 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_1_LC_9_20_4  (
            .in0(N__14947),
            .in1(N__15279),
            .in2(N__17018),
            .in3(N__14987),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(N__16892),
            .sr(N__17179));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_20_5 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_9_20_5  (
            .in0(N__21678),
            .in1(N__16981),
            .in2(_gnd_net_),
            .in3(N__20130),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(N__16892),
            .sr(N__17179));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_20_6 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_9_20_6  (
            .in0(N__15281),
            .in1(N__15365),
            .in2(N__21683),
            .in3(N__19802),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(N__16892),
            .sr(N__17179));
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_20_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_20_7 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_5_LC_9_20_7  (
            .in0(N__14983),
            .in1(N__14945),
            .in2(N__15284),
            .in3(N__19073),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(N__16892),
            .sr(N__17179));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF26P1_16_LC_9_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF26P1_16_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF26P1_16_LC_9_21_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIF26P1_16_LC_9_21_0  (
            .in0(N__20188),
            .in1(N__20259),
            .in2(N__20083),
            .in3(N__19557),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUEN44_2_LC_9_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUEN44_2_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUEN44_2_LC_9_21_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUEN44_2_LC_9_21_1  (
            .in0(N__14951),
            .in1(N__13852),
            .in2(N__13862),
            .in3(N__14771),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6L42C_31_LC_9_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6L42C_31_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6L42C_31_LC_9_21_2 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6L42C_31_LC_9_21_2  (
            .in0(N__15300),
            .in1(N__13823),
            .in2(N__13859),
            .in3(N__16974),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNI6L42C_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_RNIVV8G_0_0_LC_9_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_RNIVV8G_0_0_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.tr_state_RNIVV8G_0_0_LC_9_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.tr_state_RNIVV8G_0_0_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13853),
            .lcout(\delay_measurement_inst.N_134_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_9_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_9_21_4 .LUT_INIT=16'b0001000001010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_9_21_4  (
            .in0(N__20260),
            .in1(N__19797),
            .in2(N__15302),
            .in3(N__19558),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_160_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_9_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_9_21_5 .LUT_INIT=16'b1011101110111010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_9_21_5  (
            .in0(N__21665),
            .in1(N__16975),
            .in2(N__13856),
            .in3(N__17108),
            .lcout(\delay_measurement_inst.N_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVOI61_31_LC_9_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVOI61_31_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVOI61_31_LC_9_21_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVOI61_31_LC_9_21_6  (
            .in0(N__20898),
            .in1(N__21664),
            .in2(_gnd_net_),
            .in3(N__13851),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_reset_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_2_LC_9_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_2_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un2_startlto19_2_LC_9_21_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un2_startlto19_2_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__14787),
            .in2(_gnd_net_),
            .in3(N__14862),
            .lcout(\phase_controller_inst1.stoper_tr.un2_startlto19Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_9_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_9_22_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_9_22_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_7_LC_9_22_4  (
            .in0(N__15325),
            .in1(N__14991),
            .in2(N__19898),
            .in3(N__13793),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21120),
            .ce(),
            .sr(N__17186));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_23_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_23_3 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_9_23_3  (
            .in0(N__16985),
            .in1(N__21682),
            .in2(_gnd_net_),
            .in3(N__20189),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21115),
            .ce(N__16891),
            .sr(N__17172));
    defparam \phase_controller_inst1.start_timer_tr_LC_9_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_9_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_9_24_7 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_9_24_7  (
            .in0(N__18547),
            .in1(N__15566),
            .in2(N__21488),
            .in3(N__15210),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21110),
            .ce(),
            .sr(N__20830));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_9_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_9_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__15761),
            .in2(_gnd_net_),
            .in3(N__15189),
            .lcout(\phase_controller_inst1.N_108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_9_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_9_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_9_25_5 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \phase_controller_inst1.state_0_LC_9_25_5  (
            .in0(N__15190),
            .in1(N__15762),
            .in2(N__15245),
            .in3(N__18976),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(),
            .sr(N__20835));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_25_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_25_6  (
            .in0(N__15551),
            .in1(N__15882),
            .in2(N__15686),
            .in3(N__13961),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(),
            .sr(N__20835));
    defparam \phase_controller_slave.S1_LC_9_30_4 .C_ON=1'b0;
    defparam \phase_controller_slave.S1_LC_9_30_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S1_LC_9_30_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.S1_LC_9_30_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13937),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21100),
            .ce(),
            .sr(N__20846));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_10_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_10_9_3 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_10_9_3  (
            .in0(N__15481),
            .in1(N__15461),
            .in2(_gnd_net_),
            .in3(N__17044),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21183),
            .ce(),
            .sr(N__20760));
    defparam \delay_measurement_inst.hc_state_RNIE29G_0_LC_10_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_RNIE29G_0_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.hc_state_RNIE29G_0_LC_10_10_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \delay_measurement_inst.hc_state_RNIE29G_0_LC_10_10_0  (
            .in0(N__15419),
            .in1(N__14130),
            .in2(_gnd_net_),
            .in3(N__15432),
            .lcout(\delay_measurement_inst.N_54 ),
            .ltout(\delay_measurement_inst.N_54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_state_RNIE29G_0_0_LC_10_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_RNIE29G_0_0_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.hc_state_RNIE29G_0_0_LC_10_10_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \delay_measurement_inst.hc_state_RNIE29G_0_0_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13886),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.N_54_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_10_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_10_10_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_10_10_3  (
            .in0(N__15434),
            .in1(N__20890),
            .in2(N__14138),
            .in3(N__15421),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21177),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_10_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_10_10_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_10_10_5  (
            .in0(N__13882),
            .in1(N__20891),
            .in2(N__14171),
            .in3(N__14153),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21177),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_state_0_LC_10_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_10_10_7 .LUT_INIT=16'b0010000100110000;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_10_10_7  (
            .in0(N__15433),
            .in1(N__20889),
            .in2(N__14137),
            .in3(N__15420),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21177),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_esr_14_LC_10_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_14_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_14_LC_10_11_0 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_14_LC_10_11_0  (
            .in0(N__17833),
            .in1(N__14120),
            .in2(N__17996),
            .in3(N__17974),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21170),
            .ce(N__17681),
            .sr(N__17656));
    defparam \delay_measurement_inst.delay_hc_reg_esr_9_LC_10_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_9_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_9_LC_10_11_2 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_9_LC_10_11_2  (
            .in0(N__14210),
            .in1(N__17710),
            .in2(N__17837),
            .in3(N__14090),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21170),
            .ce(N__17681),
            .sr(N__17656));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_10_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_10_12_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_10_12_0  (
            .in0(N__14251),
            .in1(N__14063),
            .in2(N__16064),
            .in3(N__14026),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21162),
            .ce(),
            .sr(N__17657));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8R7QA_31_LC_10_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8R7QA_31_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8R7QA_31_LC_10_12_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8R7QA_31_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__14025),
            .in2(_gnd_net_),
            .in3(N__14041),
            .lcout(\delay_measurement_inst.N_54_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_10_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_10_12_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_10_12_3  (
            .in0(N__14027),
            .in1(N__14012),
            .in2(N__16102),
            .in3(N__14252),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21162),
            .ce(),
            .sr(N__17657));
    defparam \delay_measurement_inst.delay_hc_reg_ess_1_LC_10_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_ess_1_LC_10_13_0 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_ess_1_LC_10_13_0 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_ess_1_LC_10_13_0  (
            .in0(N__14258),
            .in1(N__14215),
            .in2(N__13994),
            .in3(N__14302),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21155),
            .ce(N__17682),
            .sr(N__17659));
    defparam \delay_measurement_inst.delay_hc_reg_esr_10_LC_10_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_10_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_10_LC_10_13_1 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_10_LC_10_13_1  (
            .in0(N__13976),
            .in1(N__17821),
            .in2(_gnd_net_),
            .in3(N__17708),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21155),
            .ce(N__17682),
            .sr(N__17659));
    defparam \delay_measurement_inst.delay_hc_reg_esr_4_LC_10_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_4_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_4_LC_10_13_2 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_4_LC_10_13_2  (
            .in0(N__14255),
            .in1(N__14301),
            .in2(N__14417),
            .in3(N__14222),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21155),
            .ce(N__17682),
            .sr(N__17659));
    defparam \delay_measurement_inst.delay_hc_reg_esr_18_LC_10_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_18_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_18_LC_10_13_3 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_18_LC_10_13_3  (
            .in0(N__17973),
            .in1(N__17826),
            .in2(_gnd_net_),
            .in3(N__14398),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21155),
            .ce(N__17682),
            .sr(N__17659));
    defparam \delay_measurement_inst.delay_hc_reg_esr_17_LC_10_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_17_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_17_LC_10_13_4 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_17_LC_10_13_4  (
            .in0(N__17825),
            .in1(N__14369),
            .in2(_gnd_net_),
            .in3(N__17972),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21155),
            .ce(N__17682),
            .sr(N__17659));
    defparam \delay_measurement_inst.delay_hc_reg_esr_6_LC_10_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_6_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_6_LC_10_13_5 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_6_LC_10_13_5  (
            .in0(N__14300),
            .in1(N__14257),
            .in2(N__14225),
            .in3(N__14345),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21155),
            .ce(N__17682),
            .sr(N__17659));
    defparam \delay_measurement_inst.delay_hc_reg_esr_13_LC_10_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_13_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_13_LC_10_13_6 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_13_LC_10_13_6  (
            .in0(N__17709),
            .in1(_gnd_net_),
            .in2(N__17832),
            .in3(N__14330),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21155),
            .ce(N__17682),
            .sr(N__17659));
    defparam \delay_measurement_inst.delay_hc_reg_esr_5_LC_10_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_5_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_5_LC_10_13_7 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_5_LC_10_13_7  (
            .in0(N__14299),
            .in1(N__14256),
            .in2(N__14224),
            .in3(N__14186),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21155),
            .ce(N__17682),
            .sr(N__17659));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_10_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_10_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_10_14_0 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_10_14_0  (
            .in0(N__16562),
            .in1(N__16355),
            .in2(N__17400),
            .in3(N__16682),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(N__18773),
            .sr(N__20779));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_10_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_10_14_1 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_10_14_1 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_10_14_1  (
            .in0(N__16123),
            .in1(N__16005),
            .in2(N__17242),
            .in3(N__16285),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(N__18773),
            .sr(N__20779));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_10_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_10_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_10_14_3 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_10_14_3  (
            .in0(N__16685),
            .in1(N__16565),
            .in2(N__16400),
            .in3(N__16101),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(N__18773),
            .sr(N__20779));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_14_4 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_10_14_4  (
            .in0(N__16563),
            .in1(N__16356),
            .in2(N__17363),
            .in3(N__16683),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(N__18773),
            .sr(N__20779));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_14_5 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_10_14_5  (
            .in0(N__16684),
            .in1(N__16564),
            .in2(N__16399),
            .in3(N__16063),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(N__18773),
            .sr(N__20779));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_14_6 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_14_6 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_10_14_6  (
            .in0(N__17438),
            .in1(N__17234),
            .in2(N__16011),
            .in3(N__16122),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(N__18773),
            .sr(N__20779));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_10_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_10_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_10_14_7 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_10_14_7  (
            .in0(N__16681),
            .in1(N__15973),
            .in2(N__16398),
            .in3(N__16566),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(N__18773),
            .sr(N__20779));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__14498),
            .in2(N__14492),
            .in3(N__18246),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__14483),
            .in2(N__14474),
            .in3(N__18220),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__14465),
            .in2(N__14456),
            .in3(N__18196),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__14447),
            .in2(N__14441),
            .in3(N__18163),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__14432),
            .in2(N__14426),
            .in3(N__18139),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__16814),
            .in2(N__14597),
            .in3(N__18112),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__14588),
            .in2(N__14579),
            .in3(N__18091),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__14570),
            .in2(N__14561),
            .in3(N__18064),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_16_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_16_0  (
            .in0(N__18400),
            .in1(N__16769),
            .in2(N__14552),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__16490),
            .in2(N__14543),
            .in3(N__18376),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__16808),
            .in2(N__14534),
            .in3(N__18355),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__16763),
            .in2(N__14525),
            .in3(N__19520),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__16727),
            .in2(N__14516),
            .in3(N__18331),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__16451),
            .in2(N__14507),
            .in3(N__18310),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__16298),
            .in2(N__14696),
            .in3(N__18289),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__14687),
            .in2(N__14675),
            .in3(N__18268),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__14666),
            .in2(N__14657),
            .in3(N__18478),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__14648),
            .in2(N__14639),
            .in3(N__18457),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__14630),
            .in2(N__14621),
            .in3(N__18436),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14612),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_10_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_10_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_10_18_0 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_12_LC_10_18_0  (
            .in0(N__16603),
            .in1(N__17321),
            .in2(N__16440),
            .in3(N__16713),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21131),
            .ce(N__15142),
            .sr(N__20796));
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_10_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_10_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_10_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_19_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16232),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21131),
            .ce(N__15142),
            .sr(N__20796));
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_10_18_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_10_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_10_18_2 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_11_LC_10_18_2  (
            .in0(N__16602),
            .in1(N__17282),
            .in2(N__16439),
            .in3(N__16712),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21131),
            .ce(N__15142),
            .sr(N__20796));
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_10_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_10_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_10_18_4 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_7_LC_10_18_4  (
            .in0(N__16604),
            .in1(N__16062),
            .in2(N__16441),
            .in3(N__16714),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21131),
            .ce(N__15142),
            .sr(N__20796));
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_10_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_10_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_10_18_5 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_9_LC_10_18_5  (
            .in0(N__16715),
            .in1(N__16801),
            .in2(N__17921),
            .in3(N__16428),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21131),
            .ce(N__15142),
            .sr(N__20796));
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_10_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_10_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_10_18_6 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_10_LC_10_18_6  (
            .in0(N__16601),
            .in1(N__16514),
            .in2(N__16438),
            .in3(N__16711),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21131),
            .ce(N__15142),
            .sr(N__20796));
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_10_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_10_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_10_18_7 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_15_LC_10_18_7  (
            .in0(N__17920),
            .in1(N__16415),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21131),
            .ce(N__15142),
            .sr(N__20796));
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_10_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_10_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_10_19_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_14_LC_10_19_0  (
            .in0(N__17916),
            .in1(N__16430),
            .in2(_gnd_net_),
            .in3(N__16484),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21126),
            .ce(N__15143),
            .sr(N__20802));
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_10_19_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_10_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_10_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_16_LC_10_19_1  (
            .in0(N__16265),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21126),
            .ce(N__15143),
            .sr(N__20802));
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_10_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_10_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_10_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_17_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16199),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21126),
            .ce(N__15143),
            .sr(N__20802));
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_10_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_10_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_10_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_18_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16165),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21126),
            .ce(N__15143),
            .sr(N__20802));
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_10_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_10_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_10_19_4 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_13_LC_10_19_4  (
            .in0(N__16716),
            .in1(N__16605),
            .in2(N__16756),
            .in3(N__16429),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21126),
            .ce(N__15143),
            .sr(N__20802));
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_10_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_10_20_0 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_10_20_0 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_3_LC_10_20_0  (
            .in0(N__14989),
            .in1(N__19166),
            .in2(N__15283),
            .in3(N__14950),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21122),
            .ce(N__16886),
            .sr(N__17184));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_10_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_10_20_1 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_10_20_1  (
            .in0(N__21676),
            .in1(N__20076),
            .in2(_gnd_net_),
            .in3(N__16984),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21122),
            .ce(N__16886),
            .sr(N__17184));
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_10_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_10_20_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_10_20_3 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_4_LC_10_20_3  (
            .in0(N__14949),
            .in1(N__14990),
            .in2(N__19124),
            .in3(N__15272),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21122),
            .ce(N__16886),
            .sr(N__17184));
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_10_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_10_20_4 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_2_LC_10_20_4  (
            .in0(N__14988),
            .in1(N__16999),
            .in2(N__15282),
            .in3(N__14948),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21122),
            .ce(N__16886),
            .sr(N__17184));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_10_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_10_20_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_10_20_5  (
            .in0(N__19748),
            .in1(N__21680),
            .in2(_gnd_net_),
            .in3(N__15361),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21122),
            .ce(N__16886),
            .sr(N__17184));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_10_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_10_20_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_10_20_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_10_20_6  (
            .in0(N__15362),
            .in1(N__21677),
            .in2(_gnd_net_),
            .in3(N__19702),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21122),
            .ce(N__16886),
            .sr(N__17184));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_10_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_10_20_7 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_10_20_7  (
            .in0(N__21675),
            .in1(N__19612),
            .in2(_gnd_net_),
            .in3(N__15363),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21122),
            .ce(N__16886),
            .sr(N__17184));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_2_LC_10_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_2_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_2_LC_10_21_0 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_2_LC_10_21_0  (
            .in0(N__17000),
            .in1(N__19165),
            .in2(N__19801),
            .in3(N__17114),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_21_1 .LUT_INIT=16'b1111111100110010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_10_21_1  (
            .in0(N__20257),
            .in1(N__17104),
            .in2(N__19562),
            .in3(N__16976),
            .lcout(\delay_measurement_inst.N_132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_10_21_3  (
            .in0(N__19658),
            .in1(N__19703),
            .in2(N__19613),
            .in3(N__19744),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_10_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_10_21_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_10_21_4  (
            .in0(N__17103),
            .in1(N__21666),
            .in2(_gnd_net_),
            .in3(N__20258),
            .lcout(\delay_measurement_inst.N_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_RNI5LDIC_0_LC_10_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_RNI5LDIC_0_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.tr_state_RNI5LDIC_0_LC_10_21_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \delay_measurement_inst.tr_state_RNI5LDIC_0_LC_10_21_5  (
            .in0(N__15321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17145),
            .lcout(\delay_measurement_inst.N_134_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_21_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_10_21_6  (
            .in0(N__17090),
            .in1(N__17120),
            .in2(N__19979),
            .in3(N__17084),
            .lcout(\delay_measurement_inst.N_201 ),
            .ltout(\delay_measurement_inst.N_201_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_10_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_10_21_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_10_21_7  (
            .in0(N__20256),
            .in1(_gnd_net_),
            .in2(N__15305),
            .in3(N__15301),
            .lcout(\delay_measurement_inst.N_170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_1_LC_10_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_10_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_10_22_4 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \phase_controller_inst1.state_1_LC_10_22_4  (
            .in0(N__15244),
            .in1(N__18969),
            .in2(N__19504),
            .in3(N__21227),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21112),
            .ce(),
            .sr(N__20811));
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_10_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_10_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNIR0JF_1_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__18968),
            .in2(_gnd_net_),
            .in3(N__15243),
            .lcout(\phase_controller_inst1.T01_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.T12_LC_10_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.T12_LC_10_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T12_LC_10_25_2 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \phase_controller_inst1.T12_LC_10_25_2  (
            .in0(N__15763),
            .in1(N__15214),
            .in2(N__15166),
            .in3(N__15191),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21103),
            .ce(),
            .sr(N__20826));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_10_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_10_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_10_25_3 .LUT_INIT=16'b0010000000101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_10_25_3  (
            .in0(N__15567),
            .in1(N__15889),
            .in2(N__15715),
            .in3(N__15938),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21103),
            .ce(),
            .sr(N__20826));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_10_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_10_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_10_25_6 .LUT_INIT=16'b1111000111000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_10_25_6  (
            .in0(N__15937),
            .in1(N__15488),
            .in2(N__15767),
            .in3(N__15890),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21103),
            .ce(),
            .sr(N__20826));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_10_26_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_10_26_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_10_26_4  (
            .in0(_gnd_net_),
            .in1(N__15626),
            .in2(_gnd_net_),
            .in3(N__15568),
            .lcout(\phase_controller_inst1.stoper_tr.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_9_3 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_9_3  (
            .in0(N__15482),
            .in1(N__15460),
            .in2(_gnd_net_),
            .in3(N__17040),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_181_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_prev_LC_11_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_prev_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_prev_LC_11_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.hc_prev_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15422),
            .lcout(\delay_measurement_inst.hc_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21171),
            .ce(),
            .sr(N__20761));
    defparam \delay_measurement_inst.hc_sync_1_LC_11_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_sync_1_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_sync_1_LC_11_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.hc_sync_1_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17054),
            .lcout(\delay_measurement_inst.hc_syncZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21171),
            .ce(),
            .sr(N__20761));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI84NG1_15_LC_11_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI84NG1_15_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI84NG1_15_LC_11_12_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI84NG1_15_LC_11_12_0  (
            .in0(N__15404),
            .in1(N__17797),
            .in2(_gnd_net_),
            .in3(N__18040),
            .lcout(\delay_measurement_inst.N_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_6_LC_11_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_6_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_6_LC_11_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto19_6_LC_11_12_1  (
            .in0(N__16052),
            .in1(N__16467),
            .in2(N__16097),
            .in3(N__16790),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_12_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__15389),
            .in2(_gnd_net_),
            .in3(N__20893),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21156),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_11_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_11_12_4 .LUT_INIT=16'b1010100010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto6_LC_11_12_4  (
            .in0(N__16836),
            .in1(N__17451),
            .in2(N__17408),
            .in3(N__15956),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlt8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_11_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_11_12_5 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_11_12_5  (
            .in0(N__16468),
            .in1(N__16791),
            .in2(N__16109),
            .in3(N__16028),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_11_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_11_12_6 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_11_12_6  (
            .in0(N__16789),
            .in1(N__16084),
            .in2(_gnd_net_),
            .in3(N__16051),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_11_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_11_12_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_11_12_7  (
            .in0(N__17313),
            .in1(N__17264),
            .in2(N__16031),
            .in3(N__15949),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_8_LC_11_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_8_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_8_LC_11_13_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto19_8_LC_11_13_0  (
            .in0(N__16260),
            .in1(N__16022),
            .in2(N__16194),
            .in3(N__15950),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8 ),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_start_0_LC_11_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_start_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_start_0_LC_11_13_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_start_0_LC_11_13_1  (
            .in0(N__16329),
            .in1(N__17879),
            .in2(N__15983),
            .in3(N__17217),
            .lcout(\phase_controller_inst1.stoper_hc.un3_start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_1_LC_11_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_1_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_1_LC_11_13_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto5_1_LC_11_13_2  (
            .in0(N__16283),
            .in1(N__17345),
            .in2(_gnd_net_),
            .in3(N__15972),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_2_LC_11_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_2_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_2_LC_11_13_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto19_2_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__16743),
            .in2(_gnd_net_),
            .in3(N__16506),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_4_LC_11_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_4_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_4_LC_11_13_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto19_4_LC_11_13_4  (
            .in0(N__17878),
            .in1(N__16226),
            .in2(_gnd_net_),
            .in3(N__16160),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto6_0_LC_11_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto6_0_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto6_0_LC_11_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto6_0_LC_11_13_5  (
            .in0(N__16835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16284),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_13_6  (
            .in0(N__16259),
            .in1(N__16227),
            .in2(N__16193),
            .in3(N__16161),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_LC_11_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_LC_11_13_7 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__17880),
            .in2(N__16136),
            .in3(N__16642),
            .lcout(\phase_controller_inst1.stoper_hc.un1_start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_14_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_14_0  (
            .in0(N__19302),
            .in1(N__19456),
            .in2(N__18176),
            .in3(N__21371),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21144),
            .ce(),
            .sr(N__20776));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_14_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_14_1  (
            .in0(N__21367),
            .in1(N__19305),
            .in2(N__19461),
            .in3(N__18152),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21144),
            .ce(),
            .sr(N__20776));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_14_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_14_2  (
            .in0(N__19303),
            .in1(N__19457),
            .in2(N__18128),
            .in3(N__21372),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21144),
            .ce(),
            .sr(N__20776));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_14_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_14_3  (
            .in0(N__21368),
            .in1(N__19306),
            .in2(N__19462),
            .in3(N__18101),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21144),
            .ce(),
            .sr(N__20776));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_14_4 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_14_4  (
            .in0(N__19304),
            .in1(N__19458),
            .in2(N__18080),
            .in3(N__21373),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21144),
            .ce(),
            .sr(N__20776));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_14_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_14_5  (
            .in0(N__21369),
            .in1(N__19307),
            .in2(N__19463),
            .in3(N__18053),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21144),
            .ce(),
            .sr(N__20776));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_14_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_14_6  (
            .in0(N__19301),
            .in1(N__19455),
            .in2(N__18209),
            .in3(N__21370),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21144),
            .ce(),
            .sr(N__20776));
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_15_0 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_15_0 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_15_0  (
            .in0(N__16847),
            .in1(N__16579),
            .in2(N__16412),
            .in3(N__16675),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(N__18765),
            .sr(N__20780));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_15_1 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_11_15_1  (
            .in0(N__16677),
            .in1(N__16371),
            .in2(N__16607),
            .in3(N__17278),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(N__18765),
            .sr(N__20780));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_11_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_11_15_2 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_11_15_2  (
            .in0(N__17915),
            .in1(N__16802),
            .in2(N__16414),
            .in3(N__16680),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(N__18765),
            .sr(N__20780));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_11_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_11_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_11_15_3 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_11_15_3  (
            .in0(N__16678),
            .in1(N__16372),
            .in2(N__16608),
            .in3(N__17320),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(N__18765),
            .sr(N__20780));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_15_4 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_11_15_4  (
            .in0(N__16373),
            .in1(N__16580),
            .in2(N__16757),
            .in3(N__16679),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(N__18765),
            .sr(N__20780));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_15_5 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_11_15_5  (
            .in0(N__16676),
            .in1(N__16370),
            .in2(N__16606),
            .in3(N__16513),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(N__18765),
            .sr(N__20780));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_11_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_11_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_11_15_6 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__17913),
            .in2(N__16413),
            .in3(N__16480),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(N__18765),
            .sr(N__20780));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_15_7 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_11_15_7  (
            .in0(N__17914),
            .in1(N__16366),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(N__18765),
            .sr(N__20780));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_11_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_11_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_11_16_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_11_16_0  (
            .in0(N__21249),
            .in1(N__19284),
            .in2(N__19433),
            .in3(N__21344),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21135),
            .ce(),
            .sr(N__20781));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_11_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_11_16_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_11_16_1  (
            .in0(N__21338),
            .in1(N__18248),
            .in2(_gnd_net_),
            .in3(N__21248),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_16_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_16_2  (
            .in0(N__19381),
            .in1(N__19283),
            .in2(N__16850),
            .in3(N__21343),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21135),
            .ce(),
            .sr(N__20781));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__21311),
            .in2(_gnd_net_),
            .in3(N__21246),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_11_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_11_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_11_16_4 .LUT_INIT=16'b0000010111000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_11_16_4  (
            .in0(N__21250),
            .in1(N__19285),
            .in2(N__19434),
            .in3(N__21345),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21135),
            .ce(),
            .sr(N__20781));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_11_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_11_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__21312),
            .in2(_gnd_net_),
            .in3(N__21247),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_16_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_16_6  (
            .in0(N__19281),
            .in1(N__21339),
            .in2(N__19432),
            .in3(N__18365),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21135),
            .ce(),
            .sr(N__20781));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_16_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_16_7  (
            .in0(N__19282),
            .in1(N__19382),
            .in2(N__21374),
            .in3(N__18344),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21135),
            .ce(),
            .sr(N__20781));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_17_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_17_0  (
            .in0(N__21346),
            .in1(N__19277),
            .in2(N__19435),
            .in3(N__18320),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21132),
            .ce(),
            .sr(N__20785));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_17_1 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_17_1  (
            .in0(N__19273),
            .in1(N__19392),
            .in2(N__21387),
            .in3(N__18299),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21132),
            .ce(),
            .sr(N__20785));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_17_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_17_2  (
            .in0(N__21347),
            .in1(N__19278),
            .in2(N__19436),
            .in3(N__18278),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21132),
            .ce(),
            .sr(N__20785));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_17_3 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_17_3  (
            .in0(N__19274),
            .in1(N__19393),
            .in2(N__21388),
            .in3(N__18257),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21132),
            .ce(),
            .sr(N__20785));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_17_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_17_4  (
            .in0(N__21348),
            .in1(N__19279),
            .in2(N__19437),
            .in3(N__18467),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21132),
            .ce(),
            .sr(N__20785));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_17_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_17_5  (
            .in0(N__19275),
            .in1(N__19394),
            .in2(N__21389),
            .in3(N__18446),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21132),
            .ce(),
            .sr(N__20785));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_17_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_17_6  (
            .in0(N__21349),
            .in1(N__19280),
            .in2(N__19438),
            .in3(N__18422),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21132),
            .ce(),
            .sr(N__20785));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_17_7 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_17_7  (
            .in0(N__19276),
            .in1(N__21350),
            .in2(N__18389),
            .in3(N__19407),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21132),
            .ce(),
            .sr(N__20785));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19184),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21123),
            .ce(N__21593),
            .sr(N__20797));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19142),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21123),
            .ce(N__21593),
            .sr(N__20797));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_20_5 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_20_5  (
            .in0(N__21681),
            .in1(N__16983),
            .in2(_gnd_net_),
            .in3(N__20027),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21117),
            .ce(N__16887),
            .sr(N__17183));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_11_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_11_21_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_11_21_1  (
            .in0(N__19943),
            .in1(N__20534),
            .in2(N__20570),
            .in3(N__19910),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_7_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFD841_4_LC_11_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFD841_4_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFD841_4_LC_11_21_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFD841_4_LC_11_21_2  (
            .in0(N__20131),
            .in1(N__19072),
            .in2(N__20026),
            .in3(N__19120),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_reset_i_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_11_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_11_21_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_11_21_5  (
            .in0(N__20187),
            .in1(N__20022),
            .in2(N__20084),
            .in3(N__20132),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_11_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_11_21_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_11_21_7  (
            .in0(N__20432),
            .in1(N__20465),
            .in2(N__20396),
            .in3(N__20498),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_11_22_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_11_22_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__20294),
            .in2(_gnd_net_),
            .in3(N__20342),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_0_o2_0_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_1.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17078),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_12_8_1.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_12_8_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_12_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_12_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18863),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21176),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_sync_0_LC_12_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_sync_0_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_sync_0_LC_12_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.hc_sync_0_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17060),
            .lcout(\delay_measurement_inst.hc_syncZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21169),
            .ce(),
            .sr(N__20758));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17048),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_esr_15_LC_12_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_15_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_15_LC_12_12_3 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_15_LC_12_12_3  (
            .in0(N__17820),
            .in1(N__18044),
            .in2(N__17995),
            .in3(N__17978),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21148),
            .ce(N__17690),
            .sr(N__17660));
    defparam \delay_measurement_inst.delay_hc_reg_esr_12_LC_12_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_12_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_12_LC_12_12_6 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_12_LC_12_12_6  (
            .in0(N__17717),
            .in1(N__17858),
            .in2(_gnd_net_),
            .in3(N__17819),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21148),
            .ce(N__17690),
            .sr(N__17660));
    defparam \delay_measurement_inst.delay_hc_reg_esr_11_LC_12_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_esr_11_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_esr_11_LC_12_12_7 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_esr_11_LC_12_12_7  (
            .in0(N__17818),
            .in1(N__17738),
            .in2(_gnd_net_),
            .in3(N__17716),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21148),
            .ce(N__17690),
            .sr(N__17660));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18804),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_13_4 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_13_4  (
            .in0(N__18805),
            .in1(N__18847),
            .in2(_gnd_net_),
            .in3(N__18822),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_179_i_g ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto6_LC_12_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto6_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto6_LC_12_13_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto6_LC_12_13_6  (
            .in0(N__17452),
            .in1(N__17414),
            .in2(N__17407),
            .in3(N__17355),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlt19_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_9_LC_12_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_9_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto19_9_LC_12_13_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto19_9_LC_12_13_7  (
            .in0(N__17327),
            .in1(N__17309),
            .in2(N__17285),
            .in3(N__17265),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto19Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_14_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_14_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_12_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17201),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21140),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__18247),
            .in2(N__18230),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_12_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_12_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__18221),
            .in2(_gnd_net_),
            .in3(N__18200),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_12_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__18197),
            .in2(N__18185),
            .in3(N__18167),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_12_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_12_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__18164),
            .in2(_gnd_net_),
            .in3(N__18146),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_12_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_12_15_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18143),
            .in3(N__18119),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_12_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_12_15_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18116),
            .in3(N__18095),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_12_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_12_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__18092),
            .in2(_gnd_net_),
            .in3(N__18071),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_12_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_12_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18068),
            .in3(N__18047),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_12_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_12_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__18401),
            .in2(_gnd_net_),
            .in3(N__18380),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_12_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_12_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__18377),
            .in2(_gnd_net_),
            .in3(N__18359),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_12_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_12_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__18356),
            .in2(_gnd_net_),
            .in3(N__18338),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_12_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_12_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__19519),
            .in2(_gnd_net_),
            .in3(N__18335),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_12_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_12_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__18332),
            .in2(_gnd_net_),
            .in3(N__18314),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_12_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_12_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__18311),
            .in2(_gnd_net_),
            .in3(N__18293),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_12_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_12_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__18290),
            .in2(_gnd_net_),
            .in3(N__18272),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_12_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_12_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__18269),
            .in2(_gnd_net_),
            .in3(N__18251),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_12_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_12_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__18479),
            .in2(_gnd_net_),
            .in3(N__18461),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_12_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_12_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__18458),
            .in2(_gnd_net_),
            .in3(N__18440),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_12_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_12_17_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__18437),
            .in2(_gnd_net_),
            .in3(N__18425),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_18_0  (
            .in0(N__18705),
            .in1(N__19182),
            .in2(_gnd_net_),
            .in3(N__18416),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__21121),
            .ce(N__18593),
            .sr(N__20786));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_18_1  (
            .in0(N__18700),
            .in1(N__19140),
            .in2(_gnd_net_),
            .in3(N__18413),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__21121),
            .ce(N__18593),
            .sr(N__20786));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_18_2  (
            .in0(N__18706),
            .in1(N__19092),
            .in2(_gnd_net_),
            .in3(N__18410),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__21121),
            .ce(N__18593),
            .sr(N__20786));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_18_3  (
            .in0(N__18701),
            .in1(N__19044),
            .in2(_gnd_net_),
            .in3(N__18407),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__21121),
            .ce(N__18593),
            .sr(N__20786));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_18_4  (
            .in0(N__18707),
            .in1(N__18999),
            .in2(_gnd_net_),
            .in3(N__18404),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__21121),
            .ce(N__18593),
            .sr(N__20786));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_18_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_18_5  (
            .in0(N__18702),
            .in1(N__19869),
            .in2(_gnd_net_),
            .in3(N__18506),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__21121),
            .ce(N__18593),
            .sr(N__20786));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_18_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_18_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_18_6  (
            .in0(N__18704),
            .in1(N__19821),
            .in2(_gnd_net_),
            .in3(N__18503),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__21121),
            .ce(N__18593),
            .sr(N__20786));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_18_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_18_7  (
            .in0(N__18703),
            .in1(N__19767),
            .in2(_gnd_net_),
            .in3(N__18500),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__21121),
            .ce(N__18593),
            .sr(N__20786));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_19_0  (
            .in0(N__18699),
            .in1(N__19722),
            .in2(_gnd_net_),
            .in3(N__18497),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__21116),
            .ce(N__18594),
            .sr(N__20791));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_19_1  (
            .in0(N__18711),
            .in1(N__19677),
            .in2(_gnd_net_),
            .in3(N__18494),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__21116),
            .ce(N__18594),
            .sr(N__20791));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_19_2  (
            .in0(N__18696),
            .in1(N__19632),
            .in2(_gnd_net_),
            .in3(N__18491),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__21116),
            .ce(N__18594),
            .sr(N__20791));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_19_3  (
            .in0(N__18708),
            .in1(N__19581),
            .in2(_gnd_net_),
            .in3(N__18488),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__21116),
            .ce(N__18594),
            .sr(N__20791));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_19_4  (
            .in0(N__18697),
            .in1(N__20280),
            .in2(_gnd_net_),
            .in3(N__18485),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__21116),
            .ce(N__18594),
            .sr(N__20791));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_19_5  (
            .in0(N__18709),
            .in1(N__20208),
            .in2(_gnd_net_),
            .in3(N__18482),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__21116),
            .ce(N__18594),
            .sr(N__20791));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_19_6  (
            .in0(N__18698),
            .in1(N__20151),
            .in2(_gnd_net_),
            .in3(N__18536),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__21116),
            .ce(N__18594),
            .sr(N__20791));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_19_7  (
            .in0(N__18710),
            .in1(N__20103),
            .in2(_gnd_net_),
            .in3(N__18533),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__21116),
            .ce(N__18594),
            .sr(N__20791));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_20_0  (
            .in0(N__18714),
            .in1(N__20046),
            .in2(_gnd_net_),
            .in3(N__18530),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__21111),
            .ce(N__18595),
            .sr(N__20798));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_20_1  (
            .in0(N__18718),
            .in1(N__19998),
            .in2(_gnd_net_),
            .in3(N__18527),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__21111),
            .ce(N__18595),
            .sr(N__20798));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_20_2  (
            .in0(N__18715),
            .in1(N__19962),
            .in2(_gnd_net_),
            .in3(N__18524),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__21111),
            .ce(N__18595),
            .sr(N__20798));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_20_3  (
            .in0(N__18719),
            .in1(N__19929),
            .in2(_gnd_net_),
            .in3(N__18521),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__21111),
            .ce(N__18595),
            .sr(N__20798));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_20_4  (
            .in0(N__18716),
            .in1(N__20589),
            .in2(_gnd_net_),
            .in3(N__18518),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__21111),
            .ce(N__18595),
            .sr(N__20798));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_20_5  (
            .in0(N__18720),
            .in1(N__20553),
            .in2(_gnd_net_),
            .in3(N__18515),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__21111),
            .ce(N__18595),
            .sr(N__20798));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_20_6  (
            .in0(N__18717),
            .in1(N__20517),
            .in2(_gnd_net_),
            .in3(N__18512),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__21111),
            .ce(N__18595),
            .sr(N__20798));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_20_7  (
            .in0(N__18721),
            .in1(N__20484),
            .in2(_gnd_net_),
            .in3(N__18509),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__21111),
            .ce(N__18595),
            .sr(N__20798));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_21_0  (
            .in0(N__18722),
            .in1(N__20451),
            .in2(_gnd_net_),
            .in3(N__18740),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__21107),
            .ce(N__18596),
            .sr(N__20803));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_21_1  (
            .in0(N__18712),
            .in1(N__20415),
            .in2(_gnd_net_),
            .in3(N__18737),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__21107),
            .ce(N__18596),
            .sr(N__20803));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_21_2  (
            .in0(N__18723),
            .in1(N__20376),
            .in2(_gnd_net_),
            .in3(N__18734),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__21107),
            .ce(N__18596),
            .sr(N__20803));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_21_3  (
            .in0(N__18713),
            .in1(N__20328),
            .in2(_gnd_net_),
            .in3(N__18731),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__21107),
            .ce(N__18596),
            .sr(N__20803));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_21_4  (
            .in0(N__18724),
            .in1(N__20356),
            .in2(_gnd_net_),
            .in3(N__18728),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__21107),
            .ce(N__18596),
            .sr(N__20803));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_21_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_21_5  (
            .in0(N__20308),
            .in1(N__18725),
            .in2(_gnd_net_),
            .in3(N__18599),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21107),
            .ce(N__18596),
            .sr(N__20803));
    defparam \phase_controller_inst1.state_2_LC_12_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_12_22_0 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_12_22_0  (
            .in0(N__18578),
            .in1(N__19484),
            .in2(N__18937),
            .in3(N__21226),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21104),
            .ce(),
            .sr(N__20807));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(N__18920),
            .in2(_gnd_net_),
            .in3(N__18576),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_12_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_12_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_12_24_7 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \phase_controller_inst1.state_3_LC_12_24_7  (
            .in0(N__21440),
            .in1(N__18577),
            .in2(N__18936),
            .in3(N__18554),
            .lcout(\phase_controller_inst1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21102),
            .ce(),
            .sr(N__20812));
    defparam \phase_controller_inst1.S2_LC_12_25_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_12_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_12_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_12_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18980),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21101),
            .ce(),
            .sr(N__20818));
    defparam \phase_controller_inst1.S1_LC_12_29_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_12_29_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_12_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_12_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18938),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21099),
            .ce(),
            .sr(N__20836));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20899),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC1_LC_13_8_5.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_13_8_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_13_8_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_13_8_5 (
            .in0(N__18878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21184),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_sync_0_LC_13_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_sync_0_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_sync_0_LC_13_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.tr_sync_0_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21400),
            .lcout(\delay_measurement_inst.tr_syncZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21172),
            .ce(),
            .sr(N__20759));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_13_4 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_13_13_4  (
            .in0(N__18848),
            .in1(N__18830),
            .in2(_gnd_net_),
            .in3(N__18806),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21150),
            .ce(),
            .sr(N__20762));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(N__18829),
            .in2(_gnd_net_),
            .in3(N__18803),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_178_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_1_LC_13_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_1_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_1_LC_13_15_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_1_LC_13_15_3  (
            .in0(N__19445),
            .in1(N__19238),
            .in2(_gnd_net_),
            .in3(N__21375),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_RNITN7VZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_16_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_16_5  (
            .in0(N__19239),
            .in1(N__21376),
            .in2(N__19460),
            .in3(N__19526),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21136),
            .ce(),
            .sr(N__20777));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_17_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__19500),
            .in2(_gnd_net_),
            .in3(N__21210),
            .lcout(\phase_controller_inst1.N_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__19459),
            .in2(_gnd_net_),
            .in3(N__19223),
            .lcout(\phase_controller_inst1.stoper_hc.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_13_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_18_5 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_13_18_5  (
            .in0(N__21480),
            .in1(N__19325),
            .in2(N__19272),
            .in3(N__19313),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21127),
            .ce(),
            .sr(N__20782));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__19183),
            .in2(N__19094),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__21124),
            .ce(N__21596),
            .sr(N__20787));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__19141),
            .in2(N__19046),
            .in3(N__19097),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__21124),
            .ce(N__21596),
            .sr(N__20787));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__19093),
            .in2(N__19001),
            .in3(N__19049),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__21124),
            .ce(N__21596),
            .sr(N__20787));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__19045),
            .in2(N__19871),
            .in3(N__19004),
            .lcout(\delay_measurement_inst.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__21124),
            .ce(N__21596),
            .sr(N__20787));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__19000),
            .in2(N__19823),
            .in3(N__19874),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__21124),
            .ce(N__21596),
            .sr(N__20787));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__19870),
            .in2(N__19769),
            .in3(N__19826),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__21124),
            .ce(N__21596),
            .sr(N__20787));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__19822),
            .in2(N__19724),
            .in3(N__19772),
            .lcout(\delay_measurement_inst.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__21124),
            .ce(N__21596),
            .sr(N__20787));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__19768),
            .in2(N__19679),
            .in3(N__19727),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__21124),
            .ce(N__21596),
            .sr(N__20787));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__19723),
            .in2(N__19634),
            .in3(N__19682),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__21118),
            .ce(N__21595),
            .sr(N__20792));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__19678),
            .in2(N__19583),
            .in3(N__19637),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__21118),
            .ce(N__21595),
            .sr(N__20792));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__19633),
            .in2(N__20282),
            .in3(N__19586),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__21118),
            .ce(N__21595),
            .sr(N__20792));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__19582),
            .in2(N__20210),
            .in3(N__19529),
            .lcout(\delay_measurement_inst.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__21118),
            .ce(N__21595),
            .sr(N__20792));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__20281),
            .in2(N__20153),
            .in3(N__20213),
            .lcout(\delay_measurement_inst.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__21118),
            .ce(N__21595),
            .sr(N__20792));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__20209),
            .in2(N__20105),
            .in3(N__20156),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__21118),
            .ce(N__21595),
            .sr(N__20792));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__20152),
            .in2(N__20048),
            .in3(N__20108),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__21118),
            .ce(N__21595),
            .sr(N__20792));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__20104),
            .in2(N__20000),
            .in3(N__20051),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__21118),
            .ce(N__21595),
            .sr(N__20792));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__20047),
            .in2(N__19964),
            .in3(N__20003),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__21113),
            .ce(N__21594),
            .sr(N__20799));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__19999),
            .in2(N__19931),
            .in3(N__19967),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__21113),
            .ce(N__21594),
            .sr(N__20799));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__19963),
            .in2(N__20591),
            .in3(N__19934),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__21113),
            .ce(N__21594),
            .sr(N__20799));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(N__19930),
            .in2(N__20555),
            .in3(N__19901),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__21113),
            .ce(N__21594),
            .sr(N__20799));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__20590),
            .in2(N__20519),
            .in3(N__20558),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__21113),
            .ce(N__21594),
            .sr(N__20799));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__20554),
            .in2(N__20486),
            .in3(N__20522),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__21113),
            .ce(N__21594),
            .sr(N__20799));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(N__20518),
            .in2(N__20453),
            .in3(N__20489),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__21113),
            .ce(N__21594),
            .sr(N__20799));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__20485),
            .in2(N__20417),
            .in3(N__20456),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__21113),
            .ce(N__21594),
            .sr(N__20799));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__20452),
            .in2(N__20378),
            .in3(N__20420),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__21108),
            .ce(N__21592),
            .sr(N__20804));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__20416),
            .in2(N__20330),
            .in3(N__20381),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__21108),
            .ce(N__21592),
            .sr(N__20804));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__20377),
            .in2(N__20357),
            .in3(N__20333),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__21108),
            .ce(N__21592),
            .sr(N__20804));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__20329),
            .in2(N__20309),
            .in3(N__20285),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__21108),
            .ce(N__21592),
            .sr(N__20804));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21686),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21108),
            .ce(N__21592),
            .sr(N__20804));
    defparam \phase_controller_inst1.state_4_LC_13_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_13_23_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_13_23_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__21530),
            .in2(_gnd_net_),
            .in3(N__21464),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21105),
            .ce(),
            .sr(N__20808));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_13_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_13_24_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__21554),
            .in2(_gnd_net_),
            .in3(N__21463),
            .lcout(\phase_controller_inst1.N_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR1_LC_14_8_4.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_14_8_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_14_8_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_14_8_4 (
            .in0(N__21434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21188),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR2_LC_14_9_7.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_14_9_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_14_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_14_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21422),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21185),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_14_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_14_17_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_14_17_3  (
            .in0(N__21214),
            .in1(N__21377),
            .in2(N__21263),
            .in3(N__21254),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21137),
            .ce(),
            .sr(N__20778));
endmodule // MAIN
