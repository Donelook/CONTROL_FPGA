// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 24 2025 23:36:46

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    start_stop,
    s2_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    input start_stop;
    output s2_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__48096;
    wire N__48095;
    wire N__48094;
    wire N__48085;
    wire N__48084;
    wire N__48083;
    wire N__48076;
    wire N__48075;
    wire N__48074;
    wire N__48067;
    wire N__48066;
    wire N__48065;
    wire N__48058;
    wire N__48057;
    wire N__48056;
    wire N__48049;
    wire N__48048;
    wire N__48047;
    wire N__48040;
    wire N__48039;
    wire N__48038;
    wire N__48031;
    wire N__48030;
    wire N__48029;
    wire N__48022;
    wire N__48021;
    wire N__48020;
    wire N__48013;
    wire N__48012;
    wire N__48011;
    wire N__48004;
    wire N__48003;
    wire N__48002;
    wire N__47995;
    wire N__47994;
    wire N__47993;
    wire N__47986;
    wire N__47985;
    wire N__47984;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47957;
    wire N__47954;
    wire N__47951;
    wire N__47948;
    wire N__47945;
    wire N__47940;
    wire N__47939;
    wire N__47938;
    wire N__47937;
    wire N__47936;
    wire N__47933;
    wire N__47932;
    wire N__47931;
    wire N__47930;
    wire N__47927;
    wire N__47926;
    wire N__47925;
    wire N__47924;
    wire N__47923;
    wire N__47922;
    wire N__47921;
    wire N__47918;
    wire N__47915;
    wire N__47912;
    wire N__47911;
    wire N__47910;
    wire N__47909;
    wire N__47908;
    wire N__47907;
    wire N__47906;
    wire N__47901;
    wire N__47900;
    wire N__47899;
    wire N__47896;
    wire N__47893;
    wire N__47892;
    wire N__47891;
    wire N__47886;
    wire N__47883;
    wire N__47880;
    wire N__47867;
    wire N__47854;
    wire N__47851;
    wire N__47848;
    wire N__47845;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47823;
    wire N__47820;
    wire N__47817;
    wire N__47814;
    wire N__47809;
    wire N__47804;
    wire N__47799;
    wire N__47790;
    wire N__47789;
    wire N__47786;
    wire N__47785;
    wire N__47784;
    wire N__47783;
    wire N__47782;
    wire N__47781;
    wire N__47780;
    wire N__47779;
    wire N__47778;
    wire N__47777;
    wire N__47776;
    wire N__47775;
    wire N__47774;
    wire N__47759;
    wire N__47744;
    wire N__47743;
    wire N__47742;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47734;
    wire N__47731;
    wire N__47730;
    wire N__47729;
    wire N__47726;
    wire N__47725;
    wire N__47722;
    wire N__47721;
    wire N__47716;
    wire N__47713;
    wire N__47710;
    wire N__47705;
    wire N__47702;
    wire N__47699;
    wire N__47696;
    wire N__47693;
    wire N__47688;
    wire N__47687;
    wire N__47686;
    wire N__47681;
    wire N__47676;
    wire N__47669;
    wire N__47664;
    wire N__47661;
    wire N__47658;
    wire N__47655;
    wire N__47646;
    wire N__47643;
    wire N__47640;
    wire N__47637;
    wire N__47634;
    wire N__47631;
    wire N__47630;
    wire N__47629;
    wire N__47628;
    wire N__47627;
    wire N__47626;
    wire N__47625;
    wire N__47624;
    wire N__47623;
    wire N__47622;
    wire N__47621;
    wire N__47620;
    wire N__47617;
    wire N__47616;
    wire N__47615;
    wire N__47612;
    wire N__47609;
    wire N__47606;
    wire N__47605;
    wire N__47590;
    wire N__47585;
    wire N__47574;
    wire N__47573;
    wire N__47572;
    wire N__47571;
    wire N__47570;
    wire N__47569;
    wire N__47566;
    wire N__47563;
    wire N__47558;
    wire N__47551;
    wire N__47546;
    wire N__47543;
    wire N__47542;
    wire N__47537;
    wire N__47536;
    wire N__47535;
    wire N__47532;
    wire N__47527;
    wire N__47524;
    wire N__47521;
    wire N__47518;
    wire N__47515;
    wire N__47514;
    wire N__47511;
    wire N__47506;
    wire N__47501;
    wire N__47496;
    wire N__47491;
    wire N__47488;
    wire N__47481;
    wire N__47480;
    wire N__47477;
    wire N__47474;
    wire N__47471;
    wire N__47468;
    wire N__47463;
    wire N__47462;
    wire N__47461;
    wire N__47460;
    wire N__47459;
    wire N__47458;
    wire N__47457;
    wire N__47456;
    wire N__47455;
    wire N__47454;
    wire N__47453;
    wire N__47452;
    wire N__47451;
    wire N__47450;
    wire N__47449;
    wire N__47448;
    wire N__47447;
    wire N__47446;
    wire N__47445;
    wire N__47444;
    wire N__47443;
    wire N__47442;
    wire N__47441;
    wire N__47440;
    wire N__47439;
    wire N__47438;
    wire N__47437;
    wire N__47436;
    wire N__47435;
    wire N__47434;
    wire N__47433;
    wire N__47432;
    wire N__47431;
    wire N__47430;
    wire N__47429;
    wire N__47428;
    wire N__47427;
    wire N__47426;
    wire N__47425;
    wire N__47424;
    wire N__47423;
    wire N__47422;
    wire N__47421;
    wire N__47420;
    wire N__47419;
    wire N__47418;
    wire N__47417;
    wire N__47416;
    wire N__47415;
    wire N__47414;
    wire N__47413;
    wire N__47412;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47408;
    wire N__47407;
    wire N__47406;
    wire N__47405;
    wire N__47404;
    wire N__47403;
    wire N__47402;
    wire N__47401;
    wire N__47400;
    wire N__47399;
    wire N__47398;
    wire N__47397;
    wire N__47396;
    wire N__47395;
    wire N__47394;
    wire N__47393;
    wire N__47392;
    wire N__47391;
    wire N__47390;
    wire N__47389;
    wire N__47388;
    wire N__47387;
    wire N__47386;
    wire N__47385;
    wire N__47384;
    wire N__47383;
    wire N__47382;
    wire N__47381;
    wire N__47380;
    wire N__47379;
    wire N__47378;
    wire N__47377;
    wire N__47376;
    wire N__47375;
    wire N__47374;
    wire N__47373;
    wire N__47372;
    wire N__47371;
    wire N__47370;
    wire N__47369;
    wire N__47368;
    wire N__47367;
    wire N__47366;
    wire N__47365;
    wire N__47364;
    wire N__47363;
    wire N__47362;
    wire N__47361;
    wire N__47360;
    wire N__47359;
    wire N__47358;
    wire N__47357;
    wire N__47356;
    wire N__47355;
    wire N__47354;
    wire N__47353;
    wire N__47352;
    wire N__47351;
    wire N__47350;
    wire N__47349;
    wire N__47348;
    wire N__47347;
    wire N__47346;
    wire N__47345;
    wire N__47344;
    wire N__47343;
    wire N__47342;
    wire N__47341;
    wire N__47340;
    wire N__47339;
    wire N__47338;
    wire N__47337;
    wire N__47336;
    wire N__47335;
    wire N__47334;
    wire N__47333;
    wire N__47332;
    wire N__47331;
    wire N__47330;
    wire N__47329;
    wire N__47328;
    wire N__47327;
    wire N__47326;
    wire N__47325;
    wire N__47324;
    wire N__47323;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47319;
    wire N__47318;
    wire N__47317;
    wire N__47316;
    wire N__47315;
    wire N__47314;
    wire N__47313;
    wire N__47312;
    wire N__47311;
    wire N__47310;
    wire N__47309;
    wire N__47308;
    wire N__47307;
    wire N__46992;
    wire N__46989;
    wire N__46988;
    wire N__46987;
    wire N__46986;
    wire N__46985;
    wire N__46984;
    wire N__46981;
    wire N__46978;
    wire N__46977;
    wire N__46974;
    wire N__46971;
    wire N__46968;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46946;
    wire N__46945;
    wire N__46944;
    wire N__46943;
    wire N__46942;
    wire N__46941;
    wire N__46940;
    wire N__46939;
    wire N__46938;
    wire N__46937;
    wire N__46936;
    wire N__46935;
    wire N__46934;
    wire N__46933;
    wire N__46932;
    wire N__46931;
    wire N__46930;
    wire N__46929;
    wire N__46928;
    wire N__46927;
    wire N__46926;
    wire N__46925;
    wire N__46924;
    wire N__46923;
    wire N__46922;
    wire N__46921;
    wire N__46920;
    wire N__46919;
    wire N__46918;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46913;
    wire N__46912;
    wire N__46911;
    wire N__46910;
    wire N__46909;
    wire N__46908;
    wire N__46907;
    wire N__46906;
    wire N__46905;
    wire N__46904;
    wire N__46903;
    wire N__46902;
    wire N__46901;
    wire N__46900;
    wire N__46897;
    wire N__46896;
    wire N__46895;
    wire N__46894;
    wire N__46893;
    wire N__46892;
    wire N__46891;
    wire N__46890;
    wire N__46889;
    wire N__46888;
    wire N__46887;
    wire N__46886;
    wire N__46885;
    wire N__46884;
    wire N__46883;
    wire N__46882;
    wire N__46881;
    wire N__46878;
    wire N__46877;
    wire N__46876;
    wire N__46875;
    wire N__46874;
    wire N__46873;
    wire N__46872;
    wire N__46869;
    wire N__46868;
    wire N__46867;
    wire N__46866;
    wire N__46865;
    wire N__46864;
    wire N__46863;
    wire N__46862;
    wire N__46861;
    wire N__46860;
    wire N__46859;
    wire N__46858;
    wire N__46857;
    wire N__46856;
    wire N__46855;
    wire N__46854;
    wire N__46853;
    wire N__46852;
    wire N__46851;
    wire N__46850;
    wire N__46849;
    wire N__46848;
    wire N__46847;
    wire N__46846;
    wire N__46845;
    wire N__46844;
    wire N__46843;
    wire N__46842;
    wire N__46841;
    wire N__46840;
    wire N__46837;
    wire N__46836;
    wire N__46835;
    wire N__46834;
    wire N__46833;
    wire N__46832;
    wire N__46831;
    wire N__46830;
    wire N__46829;
    wire N__46828;
    wire N__46827;
    wire N__46826;
    wire N__46825;
    wire N__46824;
    wire N__46823;
    wire N__46822;
    wire N__46821;
    wire N__46820;
    wire N__46819;
    wire N__46818;
    wire N__46817;
    wire N__46816;
    wire N__46815;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46811;
    wire N__46810;
    wire N__46809;
    wire N__46808;
    wire N__46807;
    wire N__46806;
    wire N__46805;
    wire N__46804;
    wire N__46803;
    wire N__46802;
    wire N__46521;
    wire N__46518;
    wire N__46515;
    wire N__46514;
    wire N__46511;
    wire N__46510;
    wire N__46507;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46489;
    wire N__46484;
    wire N__46481;
    wire N__46478;
    wire N__46473;
    wire N__46472;
    wire N__46471;
    wire N__46470;
    wire N__46467;
    wire N__46464;
    wire N__46461;
    wire N__46458;
    wire N__46455;
    wire N__46452;
    wire N__46447;
    wire N__46440;
    wire N__46437;
    wire N__46434;
    wire N__46433;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46422;
    wire N__46419;
    wire N__46416;
    wire N__46413;
    wire N__46410;
    wire N__46407;
    wire N__46402;
    wire N__46397;
    wire N__46394;
    wire N__46391;
    wire N__46388;
    wire N__46383;
    wire N__46382;
    wire N__46381;
    wire N__46380;
    wire N__46377;
    wire N__46374;
    wire N__46371;
    wire N__46368;
    wire N__46365;
    wire N__46362;
    wire N__46357;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46340;
    wire N__46337;
    wire N__46336;
    wire N__46333;
    wire N__46330;
    wire N__46327;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46315;
    wire N__46308;
    wire N__46307;
    wire N__46306;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46291;
    wire N__46288;
    wire N__46285;
    wire N__46280;
    wire N__46275;
    wire N__46272;
    wire N__46271;
    wire N__46268;
    wire N__46265;
    wire N__46260;
    wire N__46257;
    wire N__46256;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46248;
    wire N__46245;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46233;
    wire N__46230;
    wire N__46225;
    wire N__46222;
    wire N__46215;
    wire N__46214;
    wire N__46211;
    wire N__46208;
    wire N__46205;
    wire N__46202;
    wire N__46197;
    wire N__46194;
    wire N__46193;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46180;
    wire N__46175;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46165;
    wire N__46158;
    wire N__46157;
    wire N__46156;
    wire N__46155;
    wire N__46148;
    wire N__46147;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46135;
    wire N__46132;
    wire N__46127;
    wire N__46124;
    wire N__46121;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46107;
    wire N__46104;
    wire N__46101;
    wire N__46098;
    wire N__46097;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46070;
    wire N__46067;
    wire N__46064;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46044;
    wire N__46043;
    wire N__46040;
    wire N__46037;
    wire N__46034;
    wire N__46031;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46013;
    wire N__46010;
    wire N__46007;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45995;
    wire N__45994;
    wire N__45991;
    wire N__45988;
    wire N__45987;
    wire N__45984;
    wire N__45979;
    wire N__45976;
    wire N__45969;
    wire N__45968;
    wire N__45963;
    wire N__45960;
    wire N__45959;
    wire N__45958;
    wire N__45957;
    wire N__45956;
    wire N__45953;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45937;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45923;
    wire N__45922;
    wire N__45919;
    wire N__45916;
    wire N__45913;
    wire N__45910;
    wire N__45907;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45891;
    wire N__45890;
    wire N__45887;
    wire N__45884;
    wire N__45881;
    wire N__45878;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45863;
    wire N__45860;
    wire N__45857;
    wire N__45854;
    wire N__45851;
    wire N__45846;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45833;
    wire N__45830;
    wire N__45827;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45794;
    wire N__45791;
    wire N__45788;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45776;
    wire N__45773;
    wire N__45770;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45752;
    wire N__45751;
    wire N__45750;
    wire N__45749;
    wire N__45748;
    wire N__45745;
    wire N__45742;
    wire N__45741;
    wire N__45740;
    wire N__45739;
    wire N__45738;
    wire N__45735;
    wire N__45734;
    wire N__45733;
    wire N__45732;
    wire N__45731;
    wire N__45730;
    wire N__45727;
    wire N__45726;
    wire N__45725;
    wire N__45724;
    wire N__45723;
    wire N__45720;
    wire N__45717;
    wire N__45716;
    wire N__45715;
    wire N__45710;
    wire N__45701;
    wire N__45698;
    wire N__45691;
    wire N__45688;
    wire N__45685;
    wire N__45682;
    wire N__45675;
    wire N__45674;
    wire N__45673;
    wire N__45670;
    wire N__45661;
    wire N__45660;
    wire N__45651;
    wire N__45648;
    wire N__45641;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45609;
    wire N__45600;
    wire N__45599;
    wire N__45598;
    wire N__45597;
    wire N__45596;
    wire N__45593;
    wire N__45592;
    wire N__45591;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45583;
    wire N__45580;
    wire N__45577;
    wire N__45576;
    wire N__45575;
    wire N__45574;
    wire N__45573;
    wire N__45570;
    wire N__45569;
    wire N__45566;
    wire N__45565;
    wire N__45562;
    wire N__45561;
    wire N__45560;
    wire N__45559;
    wire N__45558;
    wire N__45553;
    wire N__45544;
    wire N__45535;
    wire N__45534;
    wire N__45533;
    wire N__45530;
    wire N__45521;
    wire N__45518;
    wire N__45517;
    wire N__45514;
    wire N__45513;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45499;
    wire N__45496;
    wire N__45495;
    wire N__45492;
    wire N__45489;
    wire N__45486;
    wire N__45473;
    wire N__45468;
    wire N__45463;
    wire N__45450;
    wire N__45449;
    wire N__45448;
    wire N__45447;
    wire N__45446;
    wire N__45445;
    wire N__45444;
    wire N__45443;
    wire N__45442;
    wire N__45441;
    wire N__45438;
    wire N__45429;
    wire N__45420;
    wire N__45419;
    wire N__45418;
    wire N__45417;
    wire N__45416;
    wire N__45415;
    wire N__45414;
    wire N__45413;
    wire N__45412;
    wire N__45411;
    wire N__45408;
    wire N__45407;
    wire N__45406;
    wire N__45405;
    wire N__45402;
    wire N__45399;
    wire N__45396;
    wire N__45383;
    wire N__45380;
    wire N__45379;
    wire N__45374;
    wire N__45371;
    wire N__45364;
    wire N__45363;
    wire N__45360;
    wire N__45353;
    wire N__45348;
    wire N__45345;
    wire N__45340;
    wire N__45337;
    wire N__45334;
    wire N__45331;
    wire N__45322;
    wire N__45315;
    wire N__45314;
    wire N__45311;
    wire N__45308;
    wire N__45305;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45282;
    wire N__45279;
    wire N__45278;
    wire N__45275;
    wire N__45272;
    wire N__45269;
    wire N__45266;
    wire N__45261;
    wire N__45258;
    wire N__45255;
    wire N__45252;
    wire N__45249;
    wire N__45248;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45222;
    wire N__45221;
    wire N__45218;
    wire N__45215;
    wire N__45210;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45192;
    wire N__45189;
    wire N__45188;
    wire N__45185;
    wire N__45182;
    wire N__45179;
    wire N__45174;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45161;
    wire N__45158;
    wire N__45155;
    wire N__45152;
    wire N__45149;
    wire N__45144;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45123;
    wire N__45120;
    wire N__45119;
    wire N__45116;
    wire N__45113;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45078;
    wire N__45077;
    wire N__45074;
    wire N__45071;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45044;
    wire N__45041;
    wire N__45038;
    wire N__45035;
    wire N__45032;
    wire N__45029;
    wire N__45026;
    wire N__45021;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45009;
    wire N__45006;
    wire N__45005;
    wire N__45002;
    wire N__44999;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44982;
    wire N__44981;
    wire N__44978;
    wire N__44975;
    wire N__44970;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44960;
    wire N__44957;
    wire N__44954;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44936;
    wire N__44933;
    wire N__44930;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44915;
    wire N__44912;
    wire N__44909;
    wire N__44904;
    wire N__44901;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44891;
    wire N__44890;
    wire N__44889;
    wire N__44888;
    wire N__44887;
    wire N__44886;
    wire N__44885;
    wire N__44884;
    wire N__44883;
    wire N__44882;
    wire N__44881;
    wire N__44880;
    wire N__44879;
    wire N__44878;
    wire N__44877;
    wire N__44876;
    wire N__44875;
    wire N__44874;
    wire N__44873;
    wire N__44868;
    wire N__44851;
    wire N__44834;
    wire N__44831;
    wire N__44828;
    wire N__44823;
    wire N__44822;
    wire N__44821;
    wire N__44820;
    wire N__44819;
    wire N__44814;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44802;
    wire N__44797;
    wire N__44794;
    wire N__44787;
    wire N__44784;
    wire N__44779;
    wire N__44772;
    wire N__44771;
    wire N__44770;
    wire N__44769;
    wire N__44768;
    wire N__44767;
    wire N__44766;
    wire N__44765;
    wire N__44764;
    wire N__44763;
    wire N__44760;
    wire N__44759;
    wire N__44758;
    wire N__44757;
    wire N__44756;
    wire N__44755;
    wire N__44754;
    wire N__44753;
    wire N__44752;
    wire N__44751;
    wire N__44750;
    wire N__44733;
    wire N__44730;
    wire N__44729;
    wire N__44726;
    wire N__44709;
    wire N__44708;
    wire N__44707;
    wire N__44702;
    wire N__44697;
    wire N__44696;
    wire N__44693;
    wire N__44690;
    wire N__44687;
    wire N__44684;
    wire N__44681;
    wire N__44676;
    wire N__44671;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44649;
    wire N__44648;
    wire N__44647;
    wire N__44644;
    wire N__44643;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44622;
    wire N__44621;
    wire N__44620;
    wire N__44615;
    wire N__44612;
    wire N__44611;
    wire N__44608;
    wire N__44607;
    wire N__44604;
    wire N__44601;
    wire N__44598;
    wire N__44595;
    wire N__44590;
    wire N__44583;
    wire N__44580;
    wire N__44577;
    wire N__44574;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44562;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44546;
    wire N__44543;
    wire N__44540;
    wire N__44535;
    wire N__44532;
    wire N__44529;
    wire N__44526;
    wire N__44525;
    wire N__44522;
    wire N__44519;
    wire N__44514;
    wire N__44511;
    wire N__44508;
    wire N__44505;
    wire N__44504;
    wire N__44501;
    wire N__44498;
    wire N__44493;
    wire N__44490;
    wire N__44487;
    wire N__44484;
    wire N__44481;
    wire N__44480;
    wire N__44477;
    wire N__44474;
    wire N__44469;
    wire N__44466;
    wire N__44463;
    wire N__44460;
    wire N__44457;
    wire N__44454;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44423;
    wire N__44420;
    wire N__44417;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44390;
    wire N__44387;
    wire N__44384;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44366;
    wire N__44363;
    wire N__44360;
    wire N__44357;
    wire N__44352;
    wire N__44349;
    wire N__44348;
    wire N__44347;
    wire N__44346;
    wire N__44345;
    wire N__44344;
    wire N__44343;
    wire N__44342;
    wire N__44341;
    wire N__44340;
    wire N__44339;
    wire N__44338;
    wire N__44337;
    wire N__44336;
    wire N__44335;
    wire N__44334;
    wire N__44333;
    wire N__44332;
    wire N__44331;
    wire N__44330;
    wire N__44329;
    wire N__44328;
    wire N__44327;
    wire N__44326;
    wire N__44325;
    wire N__44324;
    wire N__44323;
    wire N__44322;
    wire N__44321;
    wire N__44320;
    wire N__44311;
    wire N__44302;
    wire N__44293;
    wire N__44284;
    wire N__44275;
    wire N__44270;
    wire N__44261;
    wire N__44252;
    wire N__44243;
    wire N__44236;
    wire N__44229;
    wire N__44226;
    wire N__44225;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44211;
    wire N__44208;
    wire N__44207;
    wire N__44206;
    wire N__44205;
    wire N__44202;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44188;
    wire N__44183;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44156;
    wire N__44153;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44136;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44126;
    wire N__44123;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44103;
    wire N__44100;
    wire N__44099;
    wire N__44096;
    wire N__44093;
    wire N__44090;
    wire N__44087;
    wire N__44082;
    wire N__44079;
    wire N__44076;
    wire N__44073;
    wire N__44070;
    wire N__44067;
    wire N__44064;
    wire N__44063;
    wire N__44060;
    wire N__44057;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44042;
    wire N__44039;
    wire N__44036;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44018;
    wire N__44015;
    wire N__44012;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43997;
    wire N__43996;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43977;
    wire N__43974;
    wire N__43973;
    wire N__43972;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43960;
    wire N__43953;
    wire N__43950;
    wire N__43949;
    wire N__43948;
    wire N__43945;
    wire N__43942;
    wire N__43939;
    wire N__43936;
    wire N__43929;
    wire N__43926;
    wire N__43925;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43915;
    wire N__43912;
    wire N__43905;
    wire N__43902;
    wire N__43901;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43881;
    wire N__43878;
    wire N__43877;
    wire N__43876;
    wire N__43873;
    wire N__43870;
    wire N__43867;
    wire N__43864;
    wire N__43857;
    wire N__43854;
    wire N__43853;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43843;
    wire N__43840;
    wire N__43833;
    wire N__43830;
    wire N__43829;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43809;
    wire N__43806;
    wire N__43805;
    wire N__43804;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43785;
    wire N__43782;
    wire N__43781;
    wire N__43780;
    wire N__43777;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43761;
    wire N__43758;
    wire N__43757;
    wire N__43756;
    wire N__43753;
    wire N__43750;
    wire N__43747;
    wire N__43744;
    wire N__43737;
    wire N__43734;
    wire N__43733;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43713;
    wire N__43710;
    wire N__43709;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43699;
    wire N__43696;
    wire N__43689;
    wire N__43686;
    wire N__43685;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43665;
    wire N__43662;
    wire N__43661;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43648;
    wire N__43641;
    wire N__43638;
    wire N__43637;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43627;
    wire N__43624;
    wire N__43617;
    wire N__43614;
    wire N__43613;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43593;
    wire N__43590;
    wire N__43589;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43569;
    wire N__43566;
    wire N__43565;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43545;
    wire N__43542;
    wire N__43541;
    wire N__43540;
    wire N__43537;
    wire N__43534;
    wire N__43531;
    wire N__43528;
    wire N__43521;
    wire N__43518;
    wire N__43517;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43497;
    wire N__43494;
    wire N__43493;
    wire N__43492;
    wire N__43489;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43473;
    wire N__43470;
    wire N__43469;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43449;
    wire N__43446;
    wire N__43445;
    wire N__43444;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43425;
    wire N__43422;
    wire N__43421;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43385;
    wire N__43384;
    wire N__43381;
    wire N__43380;
    wire N__43377;
    wire N__43374;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43357;
    wire N__43352;
    wire N__43349;
    wire N__43344;
    wire N__43343;
    wire N__43342;
    wire N__43341;
    wire N__43340;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43332;
    wire N__43331;
    wire N__43330;
    wire N__43329;
    wire N__43328;
    wire N__43319;
    wire N__43306;
    wire N__43303;
    wire N__43302;
    wire N__43301;
    wire N__43300;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43271;
    wire N__43260;
    wire N__43259;
    wire N__43258;
    wire N__43257;
    wire N__43254;
    wire N__43253;
    wire N__43252;
    wire N__43251;
    wire N__43246;
    wire N__43243;
    wire N__43240;
    wire N__43239;
    wire N__43236;
    wire N__43235;
    wire N__43234;
    wire N__43229;
    wire N__43226;
    wire N__43221;
    wire N__43218;
    wire N__43215;
    wire N__43210;
    wire N__43207;
    wire N__43204;
    wire N__43199;
    wire N__43188;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43158;
    wire N__43157;
    wire N__43156;
    wire N__43149;
    wire N__43148;
    wire N__43145;
    wire N__43142;
    wire N__43141;
    wire N__43140;
    wire N__43139;
    wire N__43138;
    wire N__43137;
    wire N__43134;
    wire N__43131;
    wire N__43128;
    wire N__43119;
    wire N__43110;
    wire N__43109;
    wire N__43106;
    wire N__43105;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43088;
    wire N__43083;
    wire N__43080;
    wire N__43077;
    wire N__43074;
    wire N__43071;
    wire N__43068;
    wire N__43067;
    wire N__43064;
    wire N__43063;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43046;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43029;
    wire N__43026;
    wire N__43021;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43005;
    wire N__43002;
    wire N__43001;
    wire N__43000;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42969;
    wire N__42968;
    wire N__42967;
    wire N__42964;
    wire N__42961;
    wire N__42958;
    wire N__42951;
    wire N__42948;
    wire N__42947;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42930;
    wire N__42927;
    wire N__42926;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42916;
    wire N__42913;
    wire N__42906;
    wire N__42903;
    wire N__42902;
    wire N__42901;
    wire N__42898;
    wire N__42895;
    wire N__42894;
    wire N__42893;
    wire N__42890;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42873;
    wire N__42864;
    wire N__42861;
    wire N__42858;
    wire N__42857;
    wire N__42854;
    wire N__42851;
    wire N__42848;
    wire N__42845;
    wire N__42844;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42828;
    wire N__42825;
    wire N__42824;
    wire N__42823;
    wire N__42822;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42808;
    wire N__42803;
    wire N__42800;
    wire N__42799;
    wire N__42796;
    wire N__42793;
    wire N__42790;
    wire N__42783;
    wire N__42782;
    wire N__42781;
    wire N__42778;
    wire N__42777;
    wire N__42776;
    wire N__42775;
    wire N__42774;
    wire N__42773;
    wire N__42768;
    wire N__42761;
    wire N__42758;
    wire N__42753;
    wire N__42752;
    wire N__42751;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42725;
    wire N__42722;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42696;
    wire N__42693;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42680;
    wire N__42679;
    wire N__42676;
    wire N__42673;
    wire N__42670;
    wire N__42667;
    wire N__42662;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42647;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42629;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42611;
    wire N__42608;
    wire N__42607;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42584;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42506;
    wire N__42503;
    wire N__42500;
    wire N__42497;
    wire N__42494;
    wire N__42493;
    wire N__42490;
    wire N__42487;
    wire N__42484;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42276;
    wire N__42273;
    wire N__42270;
    wire N__42267;
    wire N__42264;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42231;
    wire N__42230;
    wire N__42227;
    wire N__42226;
    wire N__42225;
    wire N__42224;
    wire N__42223;
    wire N__42222;
    wire N__42221;
    wire N__42220;
    wire N__42219;
    wire N__42218;
    wire N__42217;
    wire N__42214;
    wire N__42209;
    wire N__42208;
    wire N__42207;
    wire N__42206;
    wire N__42205;
    wire N__42202;
    wire N__42199;
    wire N__42196;
    wire N__42193;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42179;
    wire N__42178;
    wire N__42177;
    wire N__42176;
    wire N__42171;
    wire N__42168;
    wire N__42151;
    wire N__42148;
    wire N__42131;
    wire N__42130;
    wire N__42129;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42106;
    wire N__42101;
    wire N__42098;
    wire N__42095;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42071;
    wire N__42068;
    wire N__42065;
    wire N__42062;
    wire N__42059;
    wire N__42056;
    wire N__42055;
    wire N__42054;
    wire N__42051;
    wire N__42048;
    wire N__42045;
    wire N__42042;
    wire N__42033;
    wire N__42030;
    wire N__42029;
    wire N__42026;
    wire N__42023;
    wire N__42020;
    wire N__42017;
    wire N__42012;
    wire N__42009;
    wire N__42008;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41998;
    wire N__41997;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41957;
    wire N__41954;
    wire N__41951;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41919;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41900;
    wire N__41899;
    wire N__41896;
    wire N__41895;
    wire N__41894;
    wire N__41893;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41881;
    wire N__41880;
    wire N__41879;
    wire N__41876;
    wire N__41873;
    wire N__41870;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41857;
    wire N__41854;
    wire N__41853;
    wire N__41852;
    wire N__41849;
    wire N__41842;
    wire N__41839;
    wire N__41836;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41812;
    wire N__41807;
    wire N__41802;
    wire N__41799;
    wire N__41798;
    wire N__41795;
    wire N__41790;
    wire N__41785;
    wire N__41780;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41765;
    wire N__41762;
    wire N__41751;
    wire N__41750;
    wire N__41749;
    wire N__41748;
    wire N__41747;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41726;
    wire N__41725;
    wire N__41722;
    wire N__41717;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41705;
    wire N__41704;
    wire N__41701;
    wire N__41698;
    wire N__41695;
    wire N__41692;
    wire N__41689;
    wire N__41686;
    wire N__41679;
    wire N__41676;
    wire N__41675;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41643;
    wire N__41640;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41619;
    wire N__41616;
    wire N__41613;
    wire N__41610;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41602;
    wire N__41599;
    wire N__41596;
    wire N__41593;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41572;
    wire N__41569;
    wire N__41566;
    wire N__41563;
    wire N__41556;
    wire N__41553;
    wire N__41550;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41533;
    wire N__41526;
    wire N__41523;
    wire N__41522;
    wire N__41519;
    wire N__41518;
    wire N__41515;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41499;
    wire N__41496;
    wire N__41493;
    wire N__41492;
    wire N__41491;
    wire N__41490;
    wire N__41487;
    wire N__41482;
    wire N__41479;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41465;
    wire N__41464;
    wire N__41463;
    wire N__41462;
    wire N__41461;
    wire N__41460;
    wire N__41457;
    wire N__41450;
    wire N__41443;
    wire N__41436;
    wire N__41433;
    wire N__41430;
    wire N__41429;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41412;
    wire N__41409;
    wire N__41406;
    wire N__41405;
    wire N__41404;
    wire N__41401;
    wire N__41396;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41367;
    wire N__41364;
    wire N__41363;
    wire N__41362;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41346;
    wire N__41343;
    wire N__41340;
    wire N__41337;
    wire N__41336;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41305;
    wire N__41302;
    wire N__41297;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41285;
    wire N__41282;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41262;
    wire N__41259;
    wire N__41258;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41239;
    wire N__41236;
    wire N__41233;
    wire N__41228;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41213;
    wire N__41212;
    wire N__41211;
    wire N__41210;
    wire N__41207;
    wire N__41200;
    wire N__41197;
    wire N__41190;
    wire N__41187;
    wire N__41186;
    wire N__41183;
    wire N__41182;
    wire N__41181;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41167;
    wire N__41164;
    wire N__41157;
    wire N__41154;
    wire N__41151;
    wire N__41150;
    wire N__41149;
    wire N__41146;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41118;
    wire N__41115;
    wire N__41114;
    wire N__41111;
    wire N__41108;
    wire N__41105;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41091;
    wire N__41090;
    wire N__41089;
    wire N__41086;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41074;
    wire N__41073;
    wire N__41072;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41058;
    wire N__41055;
    wire N__41050;
    wire N__41047;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40988;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40967;
    wire N__40964;
    wire N__40959;
    wire N__40958;
    wire N__40955;
    wire N__40954;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40940;
    wire N__40937;
    wire N__40934;
    wire N__40931;
    wire N__40928;
    wire N__40925;
    wire N__40920;
    wire N__40917;
    wire N__40916;
    wire N__40913;
    wire N__40912;
    wire N__40911;
    wire N__40908;
    wire N__40905;
    wire N__40900;
    wire N__40893;
    wire N__40890;
    wire N__40887;
    wire N__40886;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40878;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40862;
    wire N__40859;
    wire N__40854;
    wire N__40851;
    wire N__40844;
    wire N__40841;
    wire N__40836;
    wire N__40835;
    wire N__40834;
    wire N__40833;
    wire N__40832;
    wire N__40829;
    wire N__40824;
    wire N__40823;
    wire N__40822;
    wire N__40821;
    wire N__40820;
    wire N__40819;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40811;
    wire N__40810;
    wire N__40809;
    wire N__40808;
    wire N__40803;
    wire N__40802;
    wire N__40801;
    wire N__40800;
    wire N__40799;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40787;
    wire N__40786;
    wire N__40785;
    wire N__40784;
    wire N__40781;
    wire N__40778;
    wire N__40777;
    wire N__40776;
    wire N__40775;
    wire N__40770;
    wire N__40763;
    wire N__40760;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40750;
    wire N__40745;
    wire N__40744;
    wire N__40743;
    wire N__40742;
    wire N__40741;
    wire N__40740;
    wire N__40737;
    wire N__40730;
    wire N__40723;
    wire N__40716;
    wire N__40711;
    wire N__40706;
    wire N__40703;
    wire N__40700;
    wire N__40691;
    wire N__40684;
    wire N__40679;
    wire N__40674;
    wire N__40665;
    wire N__40662;
    wire N__40657;
    wire N__40644;
    wire N__40641;
    wire N__40640;
    wire N__40639;
    wire N__40636;
    wire N__40631;
    wire N__40630;
    wire N__40629;
    wire N__40628;
    wire N__40627;
    wire N__40626;
    wire N__40625;
    wire N__40624;
    wire N__40623;
    wire N__40622;
    wire N__40621;
    wire N__40620;
    wire N__40619;
    wire N__40618;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40604;
    wire N__40593;
    wire N__40590;
    wire N__40585;
    wire N__40578;
    wire N__40563;
    wire N__40562;
    wire N__40559;
    wire N__40556;
    wire N__40555;
    wire N__40554;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40541;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40519;
    wire N__40514;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40485;
    wire N__40484;
    wire N__40481;
    wire N__40478;
    wire N__40475;
    wire N__40470;
    wire N__40467;
    wire N__40464;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40454;
    wire N__40451;
    wire N__40446;
    wire N__40443;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40431;
    wire N__40428;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40416;
    wire N__40413;
    wire N__40410;
    wire N__40407;
    wire N__40404;
    wire N__40401;
    wire N__40398;
    wire N__40395;
    wire N__40392;
    wire N__40391;
    wire N__40388;
    wire N__40385;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40367;
    wire N__40364;
    wire N__40361;
    wire N__40358;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40340;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40316;
    wire N__40313;
    wire N__40310;
    wire N__40307;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40295;
    wire N__40292;
    wire N__40289;
    wire N__40286;
    wire N__40283;
    wire N__40278;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40253;
    wire N__40250;
    wire N__40247;
    wire N__40242;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40218;
    wire N__40215;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40196;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40166;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40140;
    wire N__40137;
    wire N__40134;
    wire N__40133;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40112;
    wire N__40109;
    wire N__40106;
    wire N__40103;
    wire N__40102;
    wire N__40099;
    wire N__40096;
    wire N__40093;
    wire N__40090;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40074;
    wire N__40073;
    wire N__40070;
    wire N__40067;
    wire N__40064;
    wire N__40061;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40049;
    wire N__40048;
    wire N__40047;
    wire N__40046;
    wire N__40045;
    wire N__40042;
    wire N__40037;
    wire N__40030;
    wire N__40025;
    wire N__40020;
    wire N__40019;
    wire N__40016;
    wire N__40015;
    wire N__40014;
    wire N__40011;
    wire N__40010;
    wire N__40007;
    wire N__40002;
    wire N__39999;
    wire N__39996;
    wire N__39991;
    wire N__39984;
    wire N__39981;
    wire N__39978;
    wire N__39977;
    wire N__39976;
    wire N__39973;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39952;
    wire N__39947;
    wire N__39942;
    wire N__39941;
    wire N__39940;
    wire N__39939;
    wire N__39938;
    wire N__39937;
    wire N__39936;
    wire N__39935;
    wire N__39934;
    wire N__39933;
    wire N__39932;
    wire N__39931;
    wire N__39930;
    wire N__39929;
    wire N__39928;
    wire N__39927;
    wire N__39926;
    wire N__39925;
    wire N__39924;
    wire N__39923;
    wire N__39922;
    wire N__39921;
    wire N__39920;
    wire N__39919;
    wire N__39918;
    wire N__39917;
    wire N__39908;
    wire N__39899;
    wire N__39890;
    wire N__39889;
    wire N__39888;
    wire N__39887;
    wire N__39886;
    wire N__39877;
    wire N__39868;
    wire N__39863;
    wire N__39854;
    wire N__39847;
    wire N__39838;
    wire N__39835;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39815;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39797;
    wire N__39794;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39784;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39761;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39749;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39734;
    wire N__39731;
    wire N__39728;
    wire N__39725;
    wire N__39722;
    wire N__39717;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39699;
    wire N__39698;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39675;
    wire N__39672;
    wire N__39671;
    wire N__39670;
    wire N__39669;
    wire N__39666;
    wire N__39665;
    wire N__39662;
    wire N__39657;
    wire N__39654;
    wire N__39653;
    wire N__39650;
    wire N__39647;
    wire N__39644;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39630;
    wire N__39627;
    wire N__39618;
    wire N__39615;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39603;
    wire N__39602;
    wire N__39599;
    wire N__39596;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39575;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39558;
    wire N__39555;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39534;
    wire N__39531;
    wire N__39530;
    wire N__39529;
    wire N__39528;
    wire N__39525;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39511;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39453;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39405;
    wire N__39402;
    wire N__39399;
    wire N__39396;
    wire N__39393;
    wire N__39390;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39246;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39077;
    wire N__39074;
    wire N__39071;
    wire N__39066;
    wire N__39063;
    wire N__39060;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39045;
    wire N__39042;
    wire N__39041;
    wire N__39040;
    wire N__39039;
    wire N__39038;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39030;
    wire N__39029;
    wire N__39028;
    wire N__39027;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39015;
    wire N__39010;
    wire N__39007;
    wire N__39006;
    wire N__39005;
    wire N__38998;
    wire N__38995;
    wire N__38990;
    wire N__38987;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38966;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38948;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38907;
    wire N__38904;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38892;
    wire N__38889;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38870;
    wire N__38869;
    wire N__38866;
    wire N__38863;
    wire N__38860;
    wire N__38857;
    wire N__38850;
    wire N__38847;
    wire N__38846;
    wire N__38845;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38826;
    wire N__38823;
    wire N__38822;
    wire N__38821;
    wire N__38818;
    wire N__38815;
    wire N__38812;
    wire N__38809;
    wire N__38802;
    wire N__38799;
    wire N__38798;
    wire N__38797;
    wire N__38794;
    wire N__38791;
    wire N__38788;
    wire N__38785;
    wire N__38778;
    wire N__38775;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38765;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38732;
    wire N__38731;
    wire N__38728;
    wire N__38725;
    wire N__38724;
    wire N__38721;
    wire N__38716;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38702;
    wire N__38697;
    wire N__38696;
    wire N__38695;
    wire N__38692;
    wire N__38689;
    wire N__38686;
    wire N__38683;
    wire N__38676;
    wire N__38673;
    wire N__38672;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38652;
    wire N__38649;
    wire N__38648;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38628;
    wire N__38625;
    wire N__38624;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38604;
    wire N__38601;
    wire N__38600;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38580;
    wire N__38577;
    wire N__38576;
    wire N__38575;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38556;
    wire N__38553;
    wire N__38552;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38532;
    wire N__38529;
    wire N__38528;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38508;
    wire N__38505;
    wire N__38504;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38484;
    wire N__38481;
    wire N__38480;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38460;
    wire N__38457;
    wire N__38456;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38446;
    wire N__38443;
    wire N__38436;
    wire N__38433;
    wire N__38432;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38412;
    wire N__38409;
    wire N__38408;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38388;
    wire N__38385;
    wire N__38384;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38364;
    wire N__38361;
    wire N__38360;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38340;
    wire N__38337;
    wire N__38336;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38316;
    wire N__38313;
    wire N__38312;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38282;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38265;
    wire N__38262;
    wire N__38259;
    wire N__38256;
    wire N__38255;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38238;
    wire N__38235;
    wire N__38234;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38214;
    wire N__38211;
    wire N__38210;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38190;
    wire N__38187;
    wire N__38186;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38166;
    wire N__38163;
    wire N__38162;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38142;
    wire N__38139;
    wire N__38138;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38100;
    wire N__38097;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38076;
    wire N__38075;
    wire N__38072;
    wire N__38069;
    wire N__38066;
    wire N__38063;
    wire N__38062;
    wire N__38057;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38022;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37940;
    wire N__37937;
    wire N__37936;
    wire N__37933;
    wire N__37932;
    wire N__37929;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37899;
    wire N__37894;
    wire N__37887;
    wire N__37886;
    wire N__37885;
    wire N__37884;
    wire N__37883;
    wire N__37882;
    wire N__37881;
    wire N__37876;
    wire N__37871;
    wire N__37870;
    wire N__37869;
    wire N__37866;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37853;
    wire N__37852;
    wire N__37849;
    wire N__37848;
    wire N__37845;
    wire N__37844;
    wire N__37843;
    wire N__37842;
    wire N__37841;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37810;
    wire N__37805;
    wire N__37802;
    wire N__37795;
    wire N__37790;
    wire N__37785;
    wire N__37782;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37766;
    wire N__37761;
    wire N__37752;
    wire N__37751;
    wire N__37748;
    wire N__37747;
    wire N__37744;
    wire N__37743;
    wire N__37740;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37698;
    wire N__37697;
    wire N__37696;
    wire N__37695;
    wire N__37692;
    wire N__37691;
    wire N__37690;
    wire N__37689;
    wire N__37684;
    wire N__37683;
    wire N__37682;
    wire N__37681;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37669;
    wire N__37668;
    wire N__37667;
    wire N__37666;
    wire N__37663;
    wire N__37660;
    wire N__37653;
    wire N__37652;
    wire N__37651;
    wire N__37650;
    wire N__37649;
    wire N__37648;
    wire N__37647;
    wire N__37646;
    wire N__37645;
    wire N__37642;
    wire N__37637;
    wire N__37634;
    wire N__37627;
    wire N__37624;
    wire N__37619;
    wire N__37614;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37582;
    wire N__37579;
    wire N__37566;
    wire N__37563;
    wire N__37562;
    wire N__37561;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37550;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37532;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37512;
    wire N__37511;
    wire N__37510;
    wire N__37509;
    wire N__37508;
    wire N__37499;
    wire N__37496;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37485;
    wire N__37478;
    wire N__37475;
    wire N__37474;
    wire N__37473;
    wire N__37472;
    wire N__37471;
    wire N__37470;
    wire N__37469;
    wire N__37464;
    wire N__37461;
    wire N__37452;
    wire N__37449;
    wire N__37440;
    wire N__37439;
    wire N__37438;
    wire N__37437;
    wire N__37436;
    wire N__37433;
    wire N__37430;
    wire N__37429;
    wire N__37428;
    wire N__37425;
    wire N__37424;
    wire N__37423;
    wire N__37422;
    wire N__37421;
    wire N__37418;
    wire N__37417;
    wire N__37416;
    wire N__37413;
    wire N__37412;
    wire N__37411;
    wire N__37410;
    wire N__37409;
    wire N__37402;
    wire N__37389;
    wire N__37378;
    wire N__37375;
    wire N__37374;
    wire N__37373;
    wire N__37372;
    wire N__37371;
    wire N__37368;
    wire N__37367;
    wire N__37366;
    wire N__37365;
    wire N__37362;
    wire N__37361;
    wire N__37358;
    wire N__37353;
    wire N__37350;
    wire N__37349;
    wire N__37346;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37329;
    wire N__37328;
    wire N__37325;
    wire N__37324;
    wire N__37323;
    wire N__37322;
    wire N__37321;
    wire N__37318;
    wire N__37315;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37288;
    wire N__37275;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37257;
    wire N__37242;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37234;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37224;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37196;
    wire N__37191;
    wire N__37190;
    wire N__37189;
    wire N__37188;
    wire N__37187;
    wire N__37186;
    wire N__37181;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37163;
    wire N__37162;
    wire N__37161;
    wire N__37160;
    wire N__37157;
    wire N__37156;
    wire N__37155;
    wire N__37154;
    wire N__37153;
    wire N__37150;
    wire N__37145;
    wire N__37142;
    wire N__37141;
    wire N__37138;
    wire N__37133;
    wire N__37128;
    wire N__37121;
    wire N__37118;
    wire N__37107;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37092;
    wire N__37091;
    wire N__37088;
    wire N__37083;
    wire N__37080;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37057;
    wire N__37052;
    wire N__37047;
    wire N__37046;
    wire N__37043;
    wire N__37042;
    wire N__37039;
    wire N__37038;
    wire N__37037;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__36993;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36966;
    wire N__36957;
    wire N__36956;
    wire N__36955;
    wire N__36952;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36927;
    wire N__36924;
    wire N__36915;
    wire N__36914;
    wire N__36913;
    wire N__36910;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36888;
    wire N__36885;
    wire N__36876;
    wire N__36875;
    wire N__36872;
    wire N__36871;
    wire N__36868;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36845;
    wire N__36842;
    wire N__36831;
    wire N__36828;
    wire N__36827;
    wire N__36826;
    wire N__36825;
    wire N__36824;
    wire N__36821;
    wire N__36818;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36804;
    wire N__36801;
    wire N__36792;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36784;
    wire N__36779;
    wire N__36776;
    wire N__36775;
    wire N__36774;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36753;
    wire N__36752;
    wire N__36751;
    wire N__36750;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36711;
    wire N__36702;
    wire N__36701;
    wire N__36698;
    wire N__36697;
    wire N__36694;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36683;
    wire N__36680;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36660;
    wire N__36657;
    wire N__36656;
    wire N__36655;
    wire N__36652;
    wire N__36649;
    wire N__36648;
    wire N__36645;
    wire N__36640;
    wire N__36637;
    wire N__36634;
    wire N__36631;
    wire N__36630;
    wire N__36627;
    wire N__36624;
    wire N__36621;
    wire N__36618;
    wire N__36609;
    wire N__36608;
    wire N__36607;
    wire N__36606;
    wire N__36603;
    wire N__36600;
    wire N__36597;
    wire N__36594;
    wire N__36591;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36564;
    wire N__36563;
    wire N__36562;
    wire N__36559;
    wire N__36558;
    wire N__36555;
    wire N__36552;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36540;
    wire N__36537;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36521;
    wire N__36516;
    wire N__36513;
    wire N__36512;
    wire N__36509;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36501;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36485;
    wire N__36480;
    wire N__36477;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36455;
    wire N__36454;
    wire N__36453;
    wire N__36452;
    wire N__36449;
    wire N__36448;
    wire N__36447;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36439;
    wire N__36438;
    wire N__36437;
    wire N__36436;
    wire N__36435;
    wire N__36434;
    wire N__36433;
    wire N__36432;
    wire N__36431;
    wire N__36430;
    wire N__36429;
    wire N__36416;
    wire N__36405;
    wire N__36400;
    wire N__36395;
    wire N__36392;
    wire N__36385;
    wire N__36376;
    wire N__36369;
    wire N__36366;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36348;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36318;
    wire N__36315;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36302;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36272;
    wire N__36269;
    wire N__36264;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36245;
    wire N__36244;
    wire N__36243;
    wire N__36242;
    wire N__36241;
    wire N__36240;
    wire N__36239;
    wire N__36238;
    wire N__36237;
    wire N__36236;
    wire N__36235;
    wire N__36234;
    wire N__36231;
    wire N__36230;
    wire N__36229;
    wire N__36228;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36203;
    wire N__36202;
    wire N__36201;
    wire N__36200;
    wire N__36199;
    wire N__36198;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36178;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36146;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36116;
    wire N__36105;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36048;
    wire N__36045;
    wire N__36042;
    wire N__36039;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35966;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35956;
    wire N__35951;
    wire N__35946;
    wire N__35943;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35932;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35910;
    wire N__35907;
    wire N__35906;
    wire N__35901;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35886;
    wire N__35883;
    wire N__35882;
    wire N__35879;
    wire N__35878;
    wire N__35873;
    wire N__35870;
    wire N__35867;
    wire N__35862;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35850;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35819;
    wire N__35818;
    wire N__35817;
    wire N__35814;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35798;
    wire N__35793;
    wire N__35790;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35775;
    wire N__35772;
    wire N__35769;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35754;
    wire N__35751;
    wire N__35750;
    wire N__35749;
    wire N__35746;
    wire N__35745;
    wire N__35742;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35718;
    wire N__35713;
    wire N__35706;
    wire N__35703;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35691;
    wire N__35688;
    wire N__35687;
    wire N__35684;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35670;
    wire N__35667;
    wire N__35664;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35646;
    wire N__35643;
    wire N__35640;
    wire N__35639;
    wire N__35636;
    wire N__35633;
    wire N__35628;
    wire N__35627;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35617;
    wire N__35610;
    wire N__35609;
    wire N__35608;
    wire N__35607;
    wire N__35606;
    wire N__35595;
    wire N__35592;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35580;
    wire N__35577;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35565;
    wire N__35564;
    wire N__35563;
    wire N__35562;
    wire N__35561;
    wire N__35558;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35550;
    wire N__35549;
    wire N__35544;
    wire N__35541;
    wire N__35530;
    wire N__35527;
    wire N__35522;
    wire N__35519;
    wire N__35516;
    wire N__35511;
    wire N__35510;
    wire N__35509;
    wire N__35508;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35495;
    wire N__35492;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35472;
    wire N__35467;
    wire N__35460;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35452;
    wire N__35449;
    wire N__35444;
    wire N__35439;
    wire N__35436;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35418;
    wire N__35415;
    wire N__35412;
    wire N__35411;
    wire N__35410;
    wire N__35407;
    wire N__35406;
    wire N__35403;
    wire N__35400;
    wire N__35395;
    wire N__35392;
    wire N__35385;
    wire N__35384;
    wire N__35383;
    wire N__35380;
    wire N__35377;
    wire N__35374;
    wire N__35371;
    wire N__35366;
    wire N__35361;
    wire N__35358;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35346;
    wire N__35343;
    wire N__35340;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35320;
    wire N__35313;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35298;
    wire N__35295;
    wire N__35294;
    wire N__35291;
    wire N__35290;
    wire N__35289;
    wire N__35288;
    wire N__35287;
    wire N__35286;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35256;
    wire N__35251;
    wire N__35238;
    wire N__35237;
    wire N__35232;
    wire N__35229;
    wire N__35226;
    wire N__35223;
    wire N__35222;
    wire N__35219;
    wire N__35218;
    wire N__35211;
    wire N__35208;
    wire N__35207;
    wire N__35202;
    wire N__35199;
    wire N__35198;
    wire N__35197;
    wire N__35194;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35169;
    wire N__35166;
    wire N__35165;
    wire N__35162;
    wire N__35161;
    wire N__35158;
    wire N__35157;
    wire N__35156;
    wire N__35151;
    wire N__35148;
    wire N__35143;
    wire N__35140;
    wire N__35133;
    wire N__35132;
    wire N__35129;
    wire N__35126;
    wire N__35123;
    wire N__35120;
    wire N__35119;
    wire N__35114;
    wire N__35111;
    wire N__35106;
    wire N__35103;
    wire N__35102;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35084;
    wire N__35081;
    wire N__35078;
    wire N__35073;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35065;
    wire N__35060;
    wire N__35059;
    wire N__35056;
    wire N__35055;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35009;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34993;
    wire N__34988;
    wire N__34985;
    wire N__34982;
    wire N__34979;
    wire N__34974;
    wire N__34973;
    wire N__34972;
    wire N__34971;
    wire N__34964;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34944;
    wire N__34943;
    wire N__34942;
    wire N__34941;
    wire N__34938;
    wire N__34935;
    wire N__34930;
    wire N__34927;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34878;
    wire N__34877;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34860;
    wire N__34859;
    wire N__34858;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34823;
    wire N__34820;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34793;
    wire N__34790;
    wire N__34787;
    wire N__34786;
    wire N__34785;
    wire N__34782;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34747;
    wire N__34742;
    wire N__34739;
    wire N__34734;
    wire N__34731;
    wire N__34730;
    wire N__34729;
    wire N__34726;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34690;
    wire N__34683;
    wire N__34682;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34656;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34627;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34605;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34582;
    wire N__34581;
    wire N__34580;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34563;
    wire N__34554;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34546;
    wire N__34541;
    wire N__34538;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34526;
    wire N__34523;
    wire N__34522;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34514;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34476;
    wire N__34475;
    wire N__34474;
    wire N__34473;
    wire N__34466;
    wire N__34463;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34451;
    wire N__34450;
    wire N__34449;
    wire N__34446;
    wire N__34441;
    wire N__34438;
    wire N__34431;
    wire N__34430;
    wire N__34427;
    wire N__34426;
    wire N__34423;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34415;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34395;
    wire N__34392;
    wire N__34383;
    wire N__34382;
    wire N__34381;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34369;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34357;
    wire N__34354;
    wire N__34347;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34335;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34293;
    wire N__34292;
    wire N__34291;
    wire N__34288;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34275;
    wire N__34270;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34254;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34230;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34176;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34142;
    wire N__34139;
    wire N__34136;
    wire N__34133;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34104;
    wire N__34101;
    wire N__34098;
    wire N__34095;
    wire N__34094;
    wire N__34091;
    wire N__34088;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34050;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33902;
    wire N__33901;
    wire N__33900;
    wire N__33897;
    wire N__33894;
    wire N__33889;
    wire N__33882;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33828;
    wire N__33825;
    wire N__33824;
    wire N__33821;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33804;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33768;
    wire N__33767;
    wire N__33764;
    wire N__33761;
    wire N__33756;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33743;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33730;
    wire N__33729;
    wire N__33726;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33705;
    wire N__33702;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33690;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33675;
    wire N__33674;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33645;
    wire N__33642;
    wire N__33641;
    wire N__33640;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33619;
    wire N__33616;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33584;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33572;
    wire N__33571;
    wire N__33568;
    wire N__33567;
    wire N__33558;
    wire N__33555;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33372;
    wire N__33371;
    wire N__33370;
    wire N__33369;
    wire N__33366;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33352;
    wire N__33345;
    wire N__33344;
    wire N__33343;
    wire N__33342;
    wire N__33341;
    wire N__33340;
    wire N__33339;
    wire N__33338;
    wire N__33337;
    wire N__33336;
    wire N__33335;
    wire N__33334;
    wire N__33333;
    wire N__33332;
    wire N__33323;
    wire N__33322;
    wire N__33321;
    wire N__33320;
    wire N__33319;
    wire N__33318;
    wire N__33317;
    wire N__33316;
    wire N__33315;
    wire N__33314;
    wire N__33313;
    wire N__33312;
    wire N__33311;
    wire N__33310;
    wire N__33309;
    wire N__33308;
    wire N__33307;
    wire N__33302;
    wire N__33293;
    wire N__33284;
    wire N__33281;
    wire N__33272;
    wire N__33263;
    wire N__33254;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33236;
    wire N__33221;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33155;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33141;
    wire N__33140;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33126;
    wire N__33117;
    wire N__33116;
    wire N__33115;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33103;
    wire N__33096;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33072;
    wire N__33069;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33045;
    wire N__33044;
    wire N__33041;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33011;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32949;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32924;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32874;
    wire N__32873;
    wire N__32872;
    wire N__32871;
    wire N__32870;
    wire N__32869;
    wire N__32868;
    wire N__32867;
    wire N__32866;
    wire N__32865;
    wire N__32864;
    wire N__32863;
    wire N__32862;
    wire N__32861;
    wire N__32860;
    wire N__32859;
    wire N__32858;
    wire N__32857;
    wire N__32856;
    wire N__32855;
    wire N__32840;
    wire N__32825;
    wire N__32814;
    wire N__32813;
    wire N__32812;
    wire N__32809;
    wire N__32804;
    wire N__32803;
    wire N__32800;
    wire N__32797;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32779;
    wire N__32776;
    wire N__32763;
    wire N__32762;
    wire N__32761;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32750;
    wire N__32749;
    wire N__32748;
    wire N__32747;
    wire N__32746;
    wire N__32745;
    wire N__32744;
    wire N__32743;
    wire N__32742;
    wire N__32741;
    wire N__32740;
    wire N__32739;
    wire N__32738;
    wire N__32737;
    wire N__32736;
    wire N__32735;
    wire N__32732;
    wire N__32731;
    wire N__32730;
    wire N__32729;
    wire N__32722;
    wire N__32719;
    wire N__32704;
    wire N__32689;
    wire N__32686;
    wire N__32683;
    wire N__32682;
    wire N__32679;
    wire N__32674;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32658;
    wire N__32655;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32580;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32565;
    wire N__32562;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32554;
    wire N__32549;
    wire N__32546;
    wire N__32543;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32524;
    wire N__32519;
    wire N__32516;
    wire N__32513;
    wire N__32508;
    wire N__32505;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32493;
    wire N__32492;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32478;
    wire N__32475;
    wire N__32474;
    wire N__32473;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32412;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32404;
    wire N__32403;
    wire N__32398;
    wire N__32395;
    wire N__32392;
    wire N__32389;
    wire N__32384;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32346;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32331;
    wire N__32328;
    wire N__32327;
    wire N__32324;
    wire N__32321;
    wire N__32318;
    wire N__32317;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32301;
    wire N__32298;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32290;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32274;
    wire N__32271;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32259;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32244;
    wire N__32241;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32229;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32214;
    wire N__32211;
    wire N__32210;
    wire N__32205;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32190;
    wire N__32187;
    wire N__32186;
    wire N__32185;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32169;
    wire N__32166;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32158;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32142;
    wire N__32139;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32131;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32115;
    wire N__32112;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32100;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32085;
    wire N__32082;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32074;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32058;
    wire N__32055;
    wire N__32054;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32044;
    wire N__32039;
    wire N__32034;
    wire N__32031;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32023;
    wire N__32018;
    wire N__32015;
    wire N__32012;
    wire N__32007;
    wire N__32004;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31996;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31980;
    wire N__31977;
    wire N__31976;
    wire N__31975;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31959;
    wire N__31956;
    wire N__31955;
    wire N__31950;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31928;
    wire N__31925;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31868;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31858;
    wire N__31855;
    wire N__31852;
    wire N__31849;
    wire N__31846;
    wire N__31839;
    wire N__31836;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31806;
    wire N__31803;
    wire N__31802;
    wire N__31801;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31785;
    wire N__31782;
    wire N__31781;
    wire N__31780;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31757;
    wire N__31754;
    wire N__31753;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31739;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31727;
    wire N__31724;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31709;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31697;
    wire N__31696;
    wire N__31695;
    wire N__31694;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31673;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31593;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31425;
    wire N__31422;
    wire N__31421;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31395;
    wire N__31394;
    wire N__31393;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31381;
    wire N__31374;
    wire N__31373;
    wire N__31372;
    wire N__31371;
    wire N__31368;
    wire N__31363;
    wire N__31360;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31343;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31335;
    wire N__31334;
    wire N__31333;
    wire N__31328;
    wire N__31323;
    wire N__31322;
    wire N__31317;
    wire N__31312;
    wire N__31309;
    wire N__31302;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31290;
    wire N__31287;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31275;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31190;
    wire N__31187;
    wire N__31184;
    wire N__31181;
    wire N__31178;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30887;
    wire N__30886;
    wire N__30885;
    wire N__30884;
    wire N__30883;
    wire N__30882;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30818;
    wire N__30811;
    wire N__30806;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30780;
    wire N__30777;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30708;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30683;
    wire N__30680;
    wire N__30679;
    wire N__30676;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30648;
    wire N__30647;
    wire N__30646;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30631;
    wire N__30628;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30594;
    wire N__30593;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30585;
    wire N__30582;
    wire N__30581;
    wire N__30580;
    wire N__30579;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30564;
    wire N__30561;
    wire N__30560;
    wire N__30557;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30537;
    wire N__30534;
    wire N__30525;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30501;
    wire N__30500;
    wire N__30497;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30473;
    wire N__30470;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30440;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30412;
    wire N__30409;
    wire N__30402;
    wire N__30399;
    wire N__30398;
    wire N__30395;
    wire N__30394;
    wire N__30393;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30369;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30351;
    wire N__30350;
    wire N__30347;
    wire N__30346;
    wire N__30343;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30315;
    wire N__30314;
    wire N__30313;
    wire N__30312;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30291;
    wire N__30290;
    wire N__30289;
    wire N__30286;
    wire N__30281;
    wire N__30280;
    wire N__30277;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30255;
    wire N__30254;
    wire N__30251;
    wire N__30250;
    wire N__30243;
    wire N__30240;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30203;
    wire N__30200;
    wire N__30197;
    wire N__30196;
    wire N__30189;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30171;
    wire N__30168;
    wire N__30167;
    wire N__30166;
    wire N__30159;
    wire N__30158;
    wire N__30155;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30141;
    wire N__30138;
    wire N__30137;
    wire N__30132;
    wire N__30129;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30098;
    wire N__30095;
    wire N__30094;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30072;
    wire N__30071;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30037;
    wire N__30034;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30011;
    wire N__30010;
    wire N__30003;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29978;
    wire N__29977;
    wire N__29970;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29942;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29931;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29910;
    wire N__29907;
    wire N__29904;
    wire N__29903;
    wire N__29902;
    wire N__29899;
    wire N__29894;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29861;
    wire N__29860;
    wire N__29853;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29835;
    wire N__29832;
    wire N__29831;
    wire N__29830;
    wire N__29823;
    wire N__29820;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29801;
    wire N__29800;
    wire N__29793;
    wire N__29792;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29759;
    wire N__29758;
    wire N__29755;
    wire N__29750;
    wire N__29749;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29710;
    wire N__29707;
    wire N__29702;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29676;
    wire N__29673;
    wire N__29672;
    wire N__29669;
    wire N__29668;
    wire N__29665;
    wire N__29660;
    wire N__29659;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29640;
    wire N__29637;
    wire N__29636;
    wire N__29635;
    wire N__29628;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29610;
    wire N__29607;
    wire N__29606;
    wire N__29605;
    wire N__29602;
    wire N__29599;
    wire N__29594;
    wire N__29593;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29567;
    wire N__29564;
    wire N__29563;
    wire N__29560;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29540;
    wire N__29537;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29522;
    wire N__29521;
    wire N__29518;
    wire N__29513;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29498;
    wire N__29495;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29483;
    wire N__29482;
    wire N__29477;
    wire N__29474;
    wire N__29473;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29441;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29384;
    wire N__29381;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29348;
    wire N__29345;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29285;
    wire N__29282;
    wire N__29281;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29269;
    wire N__29266;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29249;
    wire N__29248;
    wire N__29245;
    wire N__29240;
    wire N__29239;
    wire N__29234;
    wire N__29231;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29216;
    wire N__29211;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29132;
    wire N__29131;
    wire N__29126;
    wire N__29123;
    wire N__29118;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29106;
    wire N__29103;
    wire N__29102;
    wire N__29101;
    wire N__29098;
    wire N__29093;
    wire N__29088;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29055;
    wire N__29052;
    wire N__29051;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28987;
    wire N__28986;
    wire N__28983;
    wire N__28982;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28959;
    wire N__28958;
    wire N__28955;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28898;
    wire N__28897;
    wire N__28894;
    wire N__28889;
    wire N__28886;
    wire N__28883;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28869;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28854;
    wire N__28851;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28773;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28700;
    wire N__28697;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28632;
    wire N__28631;
    wire N__28630;
    wire N__28629;
    wire N__28628;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28595;
    wire N__28590;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28572;
    wire N__28571;
    wire N__28570;
    wire N__28567;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28555;
    wire N__28552;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28507;
    wire N__28504;
    wire N__28499;
    wire N__28494;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28457;
    wire N__28454;
    wire N__28453;
    wire N__28452;
    wire N__28451;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28435;
    wire N__28430;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28415;
    wire N__28414;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28399;
    wire N__28394;
    wire N__28391;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28376;
    wire N__28375;
    wire N__28368;
    wire N__28365;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28346;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28331;
    wire N__28330;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28301;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28284;
    wire N__28281;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28262;
    wire N__28261;
    wire N__28258;
    wire N__28253;
    wire N__28248;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28196;
    wire N__28195;
    wire N__28188;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28160;
    wire N__28159;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28147;
    wire N__28142;
    wire N__28139;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28094;
    wire N__28093;
    wire N__28086;
    wire N__28083;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28049;
    wire N__28048;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28032;
    wire N__28031;
    wire N__28028;
    wire N__28025;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27965;
    wire N__27964;
    wire N__27961;
    wire N__27956;
    wire N__27951;
    wire N__27948;
    wire N__27945;
    wire N__27944;
    wire N__27941;
    wire N__27940;
    wire N__27933;
    wire N__27930;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27918;
    wire N__27915;
    wire N__27914;
    wire N__27913;
    wire N__27906;
    wire N__27903;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27891;
    wire N__27888;
    wire N__27887;
    wire N__27884;
    wire N__27879;
    wire N__27876;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27864;
    wire N__27861;
    wire N__27860;
    wire N__27859;
    wire N__27858;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27842;
    wire N__27841;
    wire N__27840;
    wire N__27839;
    wire N__27838;
    wire N__27837;
    wire N__27836;
    wire N__27835;
    wire N__27834;
    wire N__27833;
    wire N__27832;
    wire N__27831;
    wire N__27830;
    wire N__27829;
    wire N__27828;
    wire N__27827;
    wire N__27826;
    wire N__27823;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27801;
    wire N__27800;
    wire N__27799;
    wire N__27798;
    wire N__27791;
    wire N__27788;
    wire N__27779;
    wire N__27778;
    wire N__27777;
    wire N__27776;
    wire N__27775;
    wire N__27774;
    wire N__27773;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27760;
    wire N__27755;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27716;
    wire N__27715;
    wire N__27714;
    wire N__27713;
    wire N__27712;
    wire N__27711;
    wire N__27710;
    wire N__27709;
    wire N__27706;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27698;
    wire N__27695;
    wire N__27686;
    wire N__27681;
    wire N__27672;
    wire N__27671;
    wire N__27670;
    wire N__27669;
    wire N__27668;
    wire N__27667;
    wire N__27666;
    wire N__27659;
    wire N__27656;
    wire N__27651;
    wire N__27644;
    wire N__27635;
    wire N__27622;
    wire N__27619;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27595;
    wire N__27592;
    wire N__27587;
    wire N__27582;
    wire N__27579;
    wire N__27574;
    wire N__27567;
    wire N__27560;
    wire N__27557;
    wire N__27556;
    wire N__27553;
    wire N__27548;
    wire N__27539;
    wire N__27536;
    wire N__27535;
    wire N__27532;
    wire N__27531;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27501;
    wire N__27496;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27467;
    wire N__27466;
    wire N__27465;
    wire N__27462;
    wire N__27457;
    wire N__27454;
    wire N__27449;
    wire N__27446;
    wire N__27441;
    wire N__27438;
    wire N__27437;
    wire N__27434;
    wire N__27433;
    wire N__27426;
    wire N__27423;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27411;
    wire N__27408;
    wire N__27407;
    wire N__27406;
    wire N__27399;
    wire N__27396;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27384;
    wire N__27381;
    wire N__27380;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27368;
    wire N__27363;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27335;
    wire N__27334;
    wire N__27327;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27309;
    wire N__27306;
    wire N__27305;
    wire N__27304;
    wire N__27297;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27239;
    wire N__27238;
    wire N__27237;
    wire N__27234;
    wire N__27233;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27225;
    wire N__27222;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27202;
    wire N__27199;
    wire N__27194;
    wire N__27189;
    wire N__27186;
    wire N__27185;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27174;
    wire N__27171;
    wire N__27166;
    wire N__27163;
    wire N__27162;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26594;
    wire N__26593;
    wire N__26592;
    wire N__26591;
    wire N__26590;
    wire N__26589;
    wire N__26588;
    wire N__26587;
    wire N__26586;
    wire N__26585;
    wire N__26584;
    wire N__26583;
    wire N__26582;
    wire N__26581;
    wire N__26580;
    wire N__26571;
    wire N__26562;
    wire N__26553;
    wire N__26544;
    wire N__26543;
    wire N__26542;
    wire N__26541;
    wire N__26540;
    wire N__26539;
    wire N__26538;
    wire N__26537;
    wire N__26536;
    wire N__26535;
    wire N__26534;
    wire N__26533;
    wire N__26532;
    wire N__26531;
    wire N__26530;
    wire N__26525;
    wire N__26520;
    wire N__26511;
    wire N__26502;
    wire N__26497;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26453;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26428;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26398;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26382;
    wire N__26379;
    wire N__26378;
    wire N__26377;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26361;
    wire N__26358;
    wire N__26357;
    wire N__26356;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26340;
    wire N__26337;
    wire N__26336;
    wire N__26333;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26318;
    wire N__26313;
    wire N__26310;
    wire N__26309;
    wire N__26306;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26291;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26265;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26257;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26220;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26212;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26189;
    wire N__26186;
    wire N__26183;
    wire N__26182;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26152;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26136;
    wire N__26133;
    wire N__26132;
    wire N__26131;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26115;
    wire N__26112;
    wire N__26111;
    wire N__26110;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26094;
    wire N__26091;
    wire N__26090;
    wire N__26087;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26077;
    wire N__26072;
    wire N__26067;
    wire N__26064;
    wire N__26063;
    wire N__26060;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26045;
    wire N__26040;
    wire N__26037;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26029;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26013;
    wire N__26010;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26002;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25986;
    wire N__25983;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25975;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25959;
    wire N__25956;
    wire N__25955;
    wire N__25950;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25935;
    wire N__25932;
    wire N__25931;
    wire N__25930;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25914;
    wire N__25911;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25899;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25884;
    wire N__25881;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25869;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25854;
    wire N__25851;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25824;
    wire N__25821;
    wire N__25820;
    wire N__25817;
    wire N__25814;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25794;
    wire N__25791;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25783;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25767;
    wire N__25764;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25756;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25713;
    wire N__25710;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25615;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25599;
    wire N__25596;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25347;
    wire N__25344;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25314;
    wire N__25311;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25266;
    wire N__25263;
    wire N__25260;
    wire N__25257;
    wire N__25254;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25227;
    wire N__25224;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25194;
    wire N__25191;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25170;
    wire N__25167;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25057;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25045;
    wire N__25040;
    wire N__25035;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25027;
    wire N__25026;
    wire N__25025;
    wire N__25024;
    wire N__25023;
    wire N__25018;
    wire N__25009;
    wire N__25006;
    wire N__25005;
    wire N__25004;
    wire N__25003;
    wire N__25002;
    wire N__25001;
    wire N__24994;
    wire N__24983;
    wire N__24982;
    wire N__24981;
    wire N__24980;
    wire N__24979;
    wire N__24978;
    wire N__24977;
    wire N__24976;
    wire N__24975;
    wire N__24974;
    wire N__24973;
    wire N__24972;
    wire N__24971;
    wire N__24970;
    wire N__24969;
    wire N__24964;
    wire N__24951;
    wire N__24950;
    wire N__24949;
    wire N__24936;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24920;
    wire N__24915;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24896;
    wire N__24895;
    wire N__24894;
    wire N__24893;
    wire N__24892;
    wire N__24891;
    wire N__24890;
    wire N__24889;
    wire N__24888;
    wire N__24887;
    wire N__24886;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24872;
    wire N__24871;
    wire N__24868;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24851;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24840;
    wire N__24829;
    wire N__24828;
    wire N__24825;
    wire N__24824;
    wire N__24823;
    wire N__24822;
    wire N__24821;
    wire N__24820;
    wire N__24819;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24804;
    wire N__24795;
    wire N__24786;
    wire N__24783;
    wire N__24782;
    wire N__24779;
    wire N__24778;
    wire N__24775;
    wire N__24770;
    wire N__24767;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24753;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24739;
    wire N__24734;
    wire N__24731;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24715;
    wire N__24702;
    wire N__24699;
    wire N__24690;
    wire N__24683;
    wire N__24672;
    wire N__24671;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24663;
    wire N__24662;
    wire N__24661;
    wire N__24660;
    wire N__24659;
    wire N__24658;
    wire N__24657;
    wire N__24656;
    wire N__24655;
    wire N__24654;
    wire N__24653;
    wire N__24652;
    wire N__24651;
    wire N__24650;
    wire N__24649;
    wire N__24648;
    wire N__24647;
    wire N__24646;
    wire N__24645;
    wire N__24642;
    wire N__24641;
    wire N__24636;
    wire N__24627;
    wire N__24624;
    wire N__24611;
    wire N__24606;
    wire N__24605;
    wire N__24604;
    wire N__24603;
    wire N__24602;
    wire N__24601;
    wire N__24588;
    wire N__24583;
    wire N__24574;
    wire N__24571;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24547;
    wire N__24540;
    wire N__24537;
    wire N__24536;
    wire N__24535;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24523;
    wire N__24518;
    wire N__24515;
    wire N__24510;
    wire N__24509;
    wire N__24508;
    wire N__24507;
    wire N__24506;
    wire N__24503;
    wire N__24502;
    wire N__24501;
    wire N__24500;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24485;
    wire N__24484;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24476;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24468;
    wire N__24467;
    wire N__24466;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24411;
    wire N__24408;
    wire N__24407;
    wire N__24404;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24336;
    wire N__24333;
    wire N__24328;
    wire N__24317;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24301;
    wire N__24298;
    wire N__24293;
    wire N__24282;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24186;
    wire N__24183;
    wire N__24180;
    wire N__24179;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24159;
    wire N__24156;
    wire N__24155;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24135;
    wire N__24132;
    wire N__24131;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24111;
    wire N__24108;
    wire N__24107;
    wire N__24106;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24087;
    wire N__24084;
    wire N__24083;
    wire N__24080;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24063;
    wire N__24060;
    wire N__24059;
    wire N__24058;
    wire N__24057;
    wire N__24048;
    wire N__24047;
    wire N__24046;
    wire N__24045;
    wire N__24044;
    wire N__24043;
    wire N__24042;
    wire N__24039;
    wire N__24034;
    wire N__24025;
    wire N__24018;
    wire N__24015;
    wire N__24014;
    wire N__24011;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23994;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23976;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23964;
    wire N__23963;
    wire N__23962;
    wire N__23961;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23944;
    wire N__23941;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23922;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23904;
    wire N__23903;
    wire N__23902;
    wire N__23899;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23889;
    wire N__23886;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23859;
    wire N__23856;
    wire N__23855;
    wire N__23854;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23823;
    wire N__23822;
    wire N__23819;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23808;
    wire N__23805;
    wire N__23800;
    wire N__23797;
    wire N__23792;
    wire N__23787;
    wire N__23784;
    wire N__23783;
    wire N__23780;
    wire N__23779;
    wire N__23776;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23657;
    wire N__23654;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23637;
    wire N__23634;
    wire N__23633;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23613;
    wire N__23610;
    wire N__23609;
    wire N__23606;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23589;
    wire N__23586;
    wire N__23585;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23288;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23280;
    wire N__23277;
    wire N__23272;
    wire N__23267;
    wire N__23262;
    wire N__23259;
    wire N__23258;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23250;
    wire N__23247;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23226;
    wire N__23225;
    wire N__23224;
    wire N__23221;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23195;
    wire N__23190;
    wire N__23189;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23150;
    wire N__23145;
    wire N__23144;
    wire N__23143;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23111;
    wire N__23106;
    wire N__23105;
    wire N__23104;
    wire N__23101;
    wire N__23100;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23079;
    wire N__23076;
    wire N__23075;
    wire N__23074;
    wire N__23073;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23051;
    wire N__23046;
    wire N__23045;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23037;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23016;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22982;
    wire N__22979;
    wire N__22978;
    wire N__22975;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22934;
    wire N__22933;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22925;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22917;
    wire N__22910;
    wire N__22901;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22846;
    wire N__22843;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22825;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22802;
    wire N__22801;
    wire N__22800;
    wire N__22797;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22736;
    wire N__22735;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22698;
    wire N__22697;
    wire N__22696;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22661;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22632;
    wire N__22631;
    wire N__22630;
    wire N__22627;
    wire N__22622;
    wire N__22617;
    wire N__22614;
    wire N__22613;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22602;
    wire N__22597;
    wire N__22592;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22565;
    wire N__22564;
    wire N__22561;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22543;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22529;
    wire N__22528;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22510;
    wire N__22507;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22490;
    wire N__22489;
    wire N__22486;
    wire N__22485;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22457;
    wire N__22456;
    wire N__22455;
    wire N__22452;
    wire N__22447;
    wire N__22444;
    wire N__22439;
    wire N__22434;
    wire N__22433;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22425;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22404;
    wire N__22403;
    wire N__22402;
    wire N__22399;
    wire N__22398;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22367;
    wire N__22366;
    wire N__22363;
    wire N__22358;
    wire N__22357;
    wire N__22352;
    wire N__22349;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22321;
    wire N__22318;
    wire N__22315;
    wire N__22314;
    wire N__22313;
    wire N__22312;
    wire N__22309;
    wire N__22304;
    wire N__22301;
    wire N__22296;
    wire N__22293;
    wire N__22284;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22273;
    wire N__22272;
    wire N__22271;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22253;
    wire N__22248;
    wire N__22245;
    wire N__22236;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22228;
    wire N__22227;
    wire N__22226;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22208;
    wire N__22201;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22191;
    wire N__22188;
    wire N__22183;
    wire N__22178;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22073;
    wire N__22072;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21746;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21722;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21698;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21683;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21582;
    wire N__21581;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21564;
    wire N__21561;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21549;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21537;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21525;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21513;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21501;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21486;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21399;
    wire N__21398;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21365;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21314;
    wire N__21311;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21296;
    wire N__21295;
    wire N__21294;
    wire N__21293;
    wire N__21292;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21284;
    wire N__21281;
    wire N__21272;
    wire N__21267;
    wire N__21266;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21254;
    wire N__21251;
    wire N__21246;
    wire N__21239;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21207;
    wire N__21206;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21194;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21182;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21170;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21155;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21129;
    wire N__21126;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21005;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20993;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20928;
    wire N__20925;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20806;
    wire N__20805;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20749;
    wire N__20744;
    wire N__20741;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20723;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20675;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20648;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20564;
    wire N__20563;
    wire N__20558;
    wire N__20555;
    wire N__20554;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20550;
    wire N__20549;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20535;
    wire N__20526;
    wire N__20517;
    wire N__20514;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20502;
    wire N__20501;
    wire N__20500;
    wire N__20499;
    wire N__20498;
    wire N__20493;
    wire N__20492;
    wire N__20491;
    wire N__20490;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20467;
    wire N__20458;
    wire N__20451;
    wire N__20448;
    wire N__20447;
    wire N__20446;
    wire N__20445;
    wire N__20444;
    wire N__20441;
    wire N__20440;
    wire N__20437;
    wire N__20436;
    wire N__20435;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20424;
    wire N__20419;
    wire N__20416;
    wire N__20409;
    wire N__20400;
    wire N__20397;
    wire N__20390;
    wire N__20387;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20300;
    wire N__20299;
    wire N__20298;
    wire N__20297;
    wire N__20296;
    wire N__20287;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20219;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20209;
    wire N__20206;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20147;
    wire N__20146;
    wire N__20141;
    wire N__20138;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20117;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20081;
    wire N__20078;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19952;
    wire N__19949;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19910;
    wire N__19909;
    wire N__19906;
    wire N__19905;
    wire N__19904;
    wire N__19901;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19893;
    wire N__19892;
    wire N__19891;
    wire N__19890;
    wire N__19887;
    wire N__19880;
    wire N__19875;
    wire N__19866;
    wire N__19865;
    wire N__19860;
    wire N__19855;
    wire N__19852;
    wire N__19845;
    wire N__19842;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19811;
    wire N__19810;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19512;
    wire N__19509;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19433;
    wire N__19432;
    wire N__19431;
    wire N__19424;
    wire N__19421;
    wire N__19420;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19404;
    wire N__19401;
    wire N__19400;
    wire N__19399;
    wire N__19398;
    wire N__19397;
    wire N__19396;
    wire N__19395;
    wire N__19392;
    wire N__19383;
    wire N__19382;
    wire N__19377;
    wire N__19376;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19353;
    wire N__19350;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19287;
    wire N__19286;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19077;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19041;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19028;
    wire N__19027;
    wire N__19026;
    wire N__19025;
    wire N__19022;
    wire N__19021;
    wire N__19018;
    wire N__19017;
    wire N__19014;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__18994;
    wire N__18991;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18966;
    wire N__18963;
    wire N__18960;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18689;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18660;
    wire N__18659;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18611;
    wire N__18606;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18594;
    wire N__18593;
    wire N__18590;
    wire N__18585;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18560;
    wire N__18559;
    wire N__18558;
    wire N__18557;
    wire N__18556;
    wire N__18555;
    wire N__18550;
    wire N__18547;
    wire N__18540;
    wire N__18537;
    wire N__18536;
    wire N__18535;
    wire N__18534;
    wire N__18533;
    wire N__18532;
    wire N__18531;
    wire N__18530;
    wire N__18529;
    wire N__18528;
    wire N__18527;
    wire N__18526;
    wire N__18525;
    wire N__18524;
    wire N__18523;
    wire N__18522;
    wire N__18521;
    wire N__18520;
    wire N__18517;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18486;
    wire N__18471;
    wire N__18466;
    wire N__18453;
    wire N__18452;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18417;
    wire N__18414;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18399;
    wire N__18396;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18381;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18363;
    wire N__18360;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18340;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18326;
    wire N__18325;
    wire N__18318;
    wire N__18315;
    wire N__18314;
    wire N__18313;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18294;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18282;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18266;
    wire N__18261;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18249;
    wire N__18248;
    wire N__18243;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.m7_2_cascade_ ;
    wire bfn_1_9_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire bfn_1_10_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire bfn_1_11_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire pwm_duty_input_7;
    wire pwm_duty_input_5;
    wire pwm_duty_input_9;
    wire pwm_duty_input_8;
    wire N_22_i_i;
    wire \current_shift_inst.PI_CTRL.m14_2 ;
    wire pwm_duty_input_10;
    wire pwm_duty_input_4;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire pwm_duty_input_0;
    wire pwm_duty_input_3;
    wire \current_shift_inst.PI_CTRL.N_19 ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_ ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire bfn_2_10_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire bfn_2_11_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire bfn_2_12_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.N_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_98 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_178 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire un7_start_stop_0_a3;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire bfn_3_8_0_;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_3_11_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_3_12_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire bfn_3_13_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire bfn_4_5_0_;
    wire un5_counter_cry_1;
    wire un5_counter_cry_2;
    wire un5_counter_cry_3;
    wire un5_counter_cry_4;
    wire un5_counter_cry_5;
    wire un5_counter_cry_6;
    wire un5_counter_cry_7;
    wire un5_counter_cry_8;
    wire bfn_4_6_0_;
    wire un5_counter_cry_9;
    wire un5_counter_cry_10;
    wire un5_counter_cry_11;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire pwm_duty_input_6;
    wire i8_mux;
    wire N_28_mux;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_4_13_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_4_14_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_4_15_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_4_16_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire counter_RNO_0Z0Z_7;
    wire counterZ0Z_7;
    wire counterZ0Z_2;
    wire counterZ0Z_1;
    wire un2_counter_5_cascade_;
    wire counterZ0Z_8;
    wire counterZ0Z_11;
    wire counterZ0Z_9;
    wire counterZ0Z_5;
    wire counterZ0Z_4;
    wire counterZ0Z_6;
    wire counterZ0Z_3;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire counter_RNO_0Z0Z_12;
    wire counterZ0Z_12;
    wire counter_RNO_0Z0Z_10;
    wire counterZ0Z_10;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire bfn_5_10_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire bfn_5_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire bfn_5_12_0_;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire bfn_5_13_0_;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire counterZ0Z_0;
    wire clk_10khz_RNIIENAZ0Z2_cascade_;
    wire clk_10khz_RNIIENAZ0Z2;
    wire un2_counter_8;
    wire un2_counter_7;
    wire un2_counter_9;
    wire clk_10khz_i;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \current_shift_inst.PI_CTRL.N_46_21_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.N_34 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.N_44 ;
    wire \current_shift_inst.PI_CTRL.N_44_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ;
    wire \current_shift_inst.PI_CTRL.N_46_21 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_2 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.N_46_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire bfn_7_19_0_;
    wire \current_shift_inst.timer_phase.counter_cry_0 ;
    wire \current_shift_inst.timer_phase.counter_cry_1 ;
    wire \current_shift_inst.timer_phase.counter_cry_2 ;
    wire \current_shift_inst.timer_phase.counter_cry_3 ;
    wire \current_shift_inst.timer_phase.counter_cry_4 ;
    wire \current_shift_inst.timer_phase.counter_cry_5 ;
    wire \current_shift_inst.timer_phase.counter_cry_6 ;
    wire \current_shift_inst.timer_phase.counter_cry_7 ;
    wire bfn_7_20_0_;
    wire \current_shift_inst.timer_phase.counter_cry_8 ;
    wire \current_shift_inst.timer_phase.counter_cry_9 ;
    wire \current_shift_inst.timer_phase.counter_cry_10 ;
    wire \current_shift_inst.timer_phase.counter_cry_11 ;
    wire \current_shift_inst.timer_phase.counter_cry_12 ;
    wire \current_shift_inst.timer_phase.counter_cry_13 ;
    wire \current_shift_inst.timer_phase.counter_cry_14 ;
    wire \current_shift_inst.timer_phase.counter_cry_15 ;
    wire bfn_7_21_0_;
    wire \current_shift_inst.timer_phase.counter_cry_16 ;
    wire \current_shift_inst.timer_phase.counter_cry_17 ;
    wire \current_shift_inst.timer_phase.counter_cry_18 ;
    wire \current_shift_inst.timer_phase.counter_cry_19 ;
    wire \current_shift_inst.timer_phase.counter_cry_20 ;
    wire \current_shift_inst.timer_phase.counter_cry_21 ;
    wire \current_shift_inst.timer_phase.counter_cry_22 ;
    wire \current_shift_inst.timer_phase.counter_cry_23 ;
    wire bfn_7_22_0_;
    wire \current_shift_inst.timer_phase.counter_cry_24 ;
    wire \current_shift_inst.timer_phase.counter_cry_25 ;
    wire \current_shift_inst.timer_phase.counter_cry_26 ;
    wire \current_shift_inst.timer_phase.counter_cry_27 ;
    wire \current_shift_inst.timer_phase.counter_cry_28 ;
    wire il_min_comp2_c;
    wire il_max_comp1_c;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_8_6_0_;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_8_7_0_;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire bfn_8_8_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire bfn_8_9_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.N_47_16 ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31 ;
    wire \current_shift_inst.PI_CTRL.N_47_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.N_76 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire N_655_g;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire bfn_8_13_0_;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire bfn_8_14_0_;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_inputZ0Z_12 ;
    wire \current_shift_inst.control_input_1_cry_11 ;
    wire \current_shift_inst.control_inputZ0Z_13 ;
    wire \current_shift_inst.control_input_1_cry_12 ;
    wire \current_shift_inst.control_inputZ0Z_14 ;
    wire \current_shift_inst.control_input_1_cry_13 ;
    wire \current_shift_inst.control_inputZ0Z_15 ;
    wire \current_shift_inst.control_input_1_cry_14 ;
    wire \current_shift_inst.control_input_1_cry_15 ;
    wire \current_shift_inst.control_inputZ0Z_16 ;
    wire bfn_8_15_0_;
    wire \current_shift_inst.control_inputZ0Z_17 ;
    wire \current_shift_inst.control_input_1_cry_16 ;
    wire \current_shift_inst.control_inputZ0Z_18 ;
    wire \current_shift_inst.control_input_1_cry_17 ;
    wire \current_shift_inst.control_inputZ0Z_19 ;
    wire \current_shift_inst.control_input_1_cry_18 ;
    wire \current_shift_inst.control_inputZ0Z_20 ;
    wire \current_shift_inst.control_input_1_cry_19 ;
    wire \current_shift_inst.control_inputZ0Z_21 ;
    wire \current_shift_inst.control_input_1_cry_20 ;
    wire \current_shift_inst.control_inputZ0Z_22 ;
    wire \current_shift_inst.control_input_1_cry_21 ;
    wire \current_shift_inst.control_inputZ0Z_23 ;
    wire \current_shift_inst.control_input_1_cry_22 ;
    wire \current_shift_inst.control_input_1_cry_23 ;
    wire \current_shift_inst.control_inputZ0Z_24 ;
    wire bfn_8_16_0_;
    wire \current_shift_inst.control_input_1_cry_24 ;
    wire bfn_8_17_0_;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_2 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_3 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_4 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_5 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_6 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_7 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_8 ;
    wire bfn_8_18_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_9 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_10 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_11 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_12 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_13 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_14 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_15 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_16 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_17 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_18 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_19 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_20 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_21 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_22 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_23 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_24 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_25 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_28 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_26 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_29 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_27 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_phase.running_i ;
    wire il_min_comp1_c;
    wire \current_shift_inst.S1_syncZ0Z0 ;
    wire \current_shift_inst.S1_syncZ0Z1 ;
    wire \current_shift_inst.S1_sync_prevZ0 ;
    wire bfn_9_13_0_;
    wire \current_shift_inst.z_i_0_31 ;
    wire \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ;
    wire \current_shift_inst.un38_control_input_0_cry_0 ;
    wire \current_shift_inst.un38_control_input_0_cry_1 ;
    wire \current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_2 ;
    wire \current_shift_inst.un38_control_input_0_cry_3 ;
    wire \current_shift_inst.un38_control_input_0_cry_4 ;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.un38_control_input_0_cry_5 ;
    wire \current_shift_inst.un38_control_input_0_cry_6 ;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire bfn_9_14_0_;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.un38_control_input_0_cry_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire \current_shift_inst.un38_control_input_0_cry_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.un38_control_input_0_cry_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.un38_control_input_0_cry_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNILORI_11 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.un38_control_input_0_cry_11 ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire \current_shift_inst.un38_control_input_0_cry_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.un38_control_input_0_cry_13 ;
    wire \current_shift_inst.un38_control_input_0_cry_14 ;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire bfn_9_15_0_;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire \current_shift_inst.un38_control_input_0_cry_15 ;
    wire \current_shift_inst.control_input_1_axb_11 ;
    wire \current_shift_inst.un38_control_input_0_cry_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ;
    wire \current_shift_inst.control_input_1_axb_12 ;
    wire \current_shift_inst.un38_control_input_0_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ;
    wire \current_shift_inst.control_input_1_axb_13 ;
    wire \current_shift_inst.un38_control_input_0_cry_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ;
    wire \current_shift_inst.control_input_1_axb_14 ;
    wire \current_shift_inst.un38_control_input_0_cry_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ;
    wire \current_shift_inst.control_input_1_axb_15 ;
    wire \current_shift_inst.un38_control_input_0_cry_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ;
    wire \current_shift_inst.control_input_1_axb_16 ;
    wire \current_shift_inst.un38_control_input_0_cry_21 ;
    wire \current_shift_inst.un38_control_input_0_cry_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ;
    wire \current_shift_inst.control_input_1_axb_17 ;
    wire bfn_9_16_0_;
    wire \current_shift_inst.control_input_1_axb_18 ;
    wire \current_shift_inst.un38_control_input_0_cry_23 ;
    wire \current_shift_inst.control_input_1_axb_19 ;
    wire \current_shift_inst.un38_control_input_0_cry_24 ;
    wire \current_shift_inst.control_input_1_axb_20 ;
    wire \current_shift_inst.un38_control_input_0_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ;
    wire \current_shift_inst.control_input_1_axb_21 ;
    wire \current_shift_inst.un38_control_input_0_cry_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ;
    wire \current_shift_inst.control_input_1_axb_22 ;
    wire \current_shift_inst.un38_control_input_0_cry_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ;
    wire \current_shift_inst.control_input_1_axb_23 ;
    wire \current_shift_inst.un38_control_input_0_cry_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ;
    wire \current_shift_inst.control_input_1_axb_24 ;
    wire \current_shift_inst.un38_control_input_0_cry_29 ;
    wire \current_shift_inst.un38_control_input_0_cry_30 ;
    wire \current_shift_inst.control_input_1_cry_24_THRU_CO ;
    wire bfn_9_17_0_;
    wire \current_shift_inst.control_inputZ0Z_25 ;
    wire \current_shift_inst.phase_valid_RNISLORZ0Z2 ;
    wire bfn_9_18_0_;
    wire \current_shift_inst.z_5_cry_1 ;
    wire \current_shift_inst.z_5_cry_2 ;
    wire \current_shift_inst.z_5_cry_3 ;
    wire \current_shift_inst.z_5_cry_4 ;
    wire \current_shift_inst.z_5_cry_5 ;
    wire \current_shift_inst.z_5_cry_6 ;
    wire \current_shift_inst.z_5_cry_7 ;
    wire \current_shift_inst.z_5_cry_8 ;
    wire \current_shift_inst.elapsed_time_ns_phase_9 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.elapsed_time_ns_phase_10 ;
    wire \current_shift_inst.z_5_cry_9 ;
    wire \current_shift_inst.z_5_cry_10 ;
    wire \current_shift_inst.z_5_cry_11 ;
    wire \current_shift_inst.z_5_cry_12 ;
    wire \current_shift_inst.z_5_cry_13 ;
    wire \current_shift_inst.z_5_cry_14 ;
    wire \current_shift_inst.z_5_cry_15 ;
    wire \current_shift_inst.z_5_cry_16 ;
    wire bfn_9_20_0_;
    wire \current_shift_inst.elapsed_time_ns_phase_18 ;
    wire \current_shift_inst.z_5_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_phase_19 ;
    wire \current_shift_inst.z_5_cry_18 ;
    wire \current_shift_inst.elapsed_time_ns_phase_20 ;
    wire \current_shift_inst.z_5_cry_19 ;
    wire \current_shift_inst.elapsed_time_ns_phase_21 ;
    wire \current_shift_inst.z_5_cry_20 ;
    wire \current_shift_inst.z_5_cry_21 ;
    wire \current_shift_inst.z_5_cry_22 ;
    wire \current_shift_inst.z_5_cry_23 ;
    wire \current_shift_inst.z_5_cry_24 ;
    wire bfn_9_21_0_;
    wire \current_shift_inst.z_5_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_phase_27 ;
    wire \current_shift_inst.z_5_cry_26 ;
    wire \current_shift_inst.elapsed_time_ns_phase_28 ;
    wire \current_shift_inst.z_5_cry_27 ;
    wire \current_shift_inst.elapsed_time_ns_phase_29 ;
    wire \current_shift_inst.z_5_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.z_5_cry_29 ;
    wire \current_shift_inst.z_5_cry_30 ;
    wire il_min_comp2_D1;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_5_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_ ;
    wire il_min_comp1_D1;
    wire measured_delay_hc_22;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ;
    wire \current_shift_inst.elapsed_time_ns_phase_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ;
    wire \current_shift_inst.elapsed_time_ns_phase_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ;
    wire \current_shift_inst.elapsed_time_ns_phase_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ;
    wire \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI190J_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ;
    wire \current_shift_inst.elapsed_time_ns_phase_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ;
    wire \current_shift_inst.elapsed_time_ns_phase_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ;
    wire \current_shift_inst.elapsed_time_ns_phase_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ;
    wire \current_shift_inst.elapsed_time_ns_phase_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ;
    wire \current_shift_inst.elapsed_time_ns_phase_12 ;
    wire \current_shift_inst.elapsed_time_ns_phase_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ;
    wire \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_1 ;
    wire \current_shift_inst.N_1633_i ;
    wire \current_shift_inst.timer_phase.counterZ0Z_0 ;
    wire \current_shift_inst.timer_phase.N_188_i_g ;
    wire \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_3 ;
    wire \current_shift_inst.elapsed_time_ns_phase_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_ ;
    wire \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_4 ;
    wire \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ;
    wire G_406;
    wire bfn_10_17_0_;
    wire \current_shift_inst.elapsed_time_ns_phase_1 ;
    wire G_405;
    wire \current_shift_inst.z_cry_0 ;
    wire \current_shift_inst.z_5_2 ;
    wire \current_shift_inst.z_cry_1 ;
    wire \current_shift_inst.z_5_3 ;
    wire \current_shift_inst.z_cry_2 ;
    wire \current_shift_inst.z_5_4 ;
    wire \current_shift_inst.z_cry_3 ;
    wire \current_shift_inst.z_5_5 ;
    wire \current_shift_inst.z_cry_4 ;
    wire \current_shift_inst.z_5_6 ;
    wire \current_shift_inst.z_cry_5 ;
    wire \current_shift_inst.z_5_7 ;
    wire \current_shift_inst.z_cry_6 ;
    wire \current_shift_inst.z_cry_7 ;
    wire \current_shift_inst.z_5_8 ;
    wire bfn_10_18_0_;
    wire \current_shift_inst.z_5_9 ;
    wire \current_shift_inst.z_cry_8 ;
    wire \current_shift_inst.z_5_10 ;
    wire \current_shift_inst.z_cry_9 ;
    wire \current_shift_inst.z_5_11 ;
    wire \current_shift_inst.z_cry_10 ;
    wire \current_shift_inst.z_5_12 ;
    wire \current_shift_inst.z_cry_11 ;
    wire \current_shift_inst.z_5_13 ;
    wire \current_shift_inst.z_cry_12 ;
    wire \current_shift_inst.z_5_14 ;
    wire \current_shift_inst.z_cry_13 ;
    wire \current_shift_inst.z_5_15 ;
    wire \current_shift_inst.z_cry_14 ;
    wire \current_shift_inst.z_cry_15 ;
    wire \current_shift_inst.z_5_16 ;
    wire bfn_10_19_0_;
    wire \current_shift_inst.z_5_17 ;
    wire \current_shift_inst.z_cry_16 ;
    wire \current_shift_inst.z_5_18 ;
    wire \current_shift_inst.z_cry_17 ;
    wire \current_shift_inst.z_5_19 ;
    wire \current_shift_inst.z_cry_18 ;
    wire \current_shift_inst.z_5_20 ;
    wire \current_shift_inst.z_cry_19 ;
    wire \current_shift_inst.z_5_21 ;
    wire \current_shift_inst.z_cry_20 ;
    wire \current_shift_inst.z_5_22 ;
    wire \current_shift_inst.z_cry_21 ;
    wire \current_shift_inst.z_5_23 ;
    wire \current_shift_inst.z_cry_22 ;
    wire \current_shift_inst.z_cry_23 ;
    wire \current_shift_inst.z_5_24 ;
    wire bfn_10_20_0_;
    wire \current_shift_inst.z_5_25 ;
    wire \current_shift_inst.z_cry_24 ;
    wire \current_shift_inst.z_5_26 ;
    wire \current_shift_inst.z_cry_25 ;
    wire \current_shift_inst.z_5_27 ;
    wire \current_shift_inst.z_cry_26 ;
    wire \current_shift_inst.z_5_28 ;
    wire \current_shift_inst.z_cry_27 ;
    wire \current_shift_inst.z_5_29 ;
    wire \current_shift_inst.z_cry_28 ;
    wire \current_shift_inst.z_5_30 ;
    wire \current_shift_inst.z_cry_29 ;
    wire \current_shift_inst.z_5_cry_30_THRU_CO ;
    wire \current_shift_inst.z_cry_30 ;
    wire measured_delay_hc_21;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0_cascade_ ;
    wire measured_delay_hc_20;
    wire measured_delay_hc_23;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlt30_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_6 ;
    wire \current_shift_inst.timer_s1.N_187_i ;
    wire \current_shift_inst.phase_validZ0 ;
    wire measured_delay_hc_27;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ;
    wire \current_shift_inst.elapsed_time_ns_phase_6 ;
    wire \current_shift_inst.elapsed_time_ns_phase_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un4_control_input_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_1_fast_31 ;
    wire \current_shift_inst.un38_control_input_0 ;
    wire bfn_11_16_0_;
    wire \current_shift_inst.un4_control_input_axb_2 ;
    wire \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_1 ;
    wire \current_shift_inst.un4_control_input_axb_3 ;
    wire \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_2 ;
    wire \current_shift_inst.un4_control_input_axb_4 ;
    wire \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_3 ;
    wire \current_shift_inst.un4_control_input_axb_5 ;
    wire \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_4 ;
    wire \current_shift_inst.un4_control_input_axb_6 ;
    wire \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_5 ;
    wire \current_shift_inst.un4_control_input_axb_7 ;
    wire \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_6 ;
    wire \current_shift_inst.un4_control_input_axb_8 ;
    wire \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_7 ;
    wire \current_shift_inst.un4_control_input_cry_8 ;
    wire \current_shift_inst.un4_control_input_axb_9 ;
    wire \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ;
    wire bfn_11_17_0_;
    wire \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ;
    wire \current_shift_inst.un4_control_input_cry_9 ;
    wire \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ;
    wire \current_shift_inst.un4_control_input_cry_10 ;
    wire \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ;
    wire \current_shift_inst.un4_control_input_cry_11 ;
    wire \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ;
    wire \current_shift_inst.un4_control_input_cry_12 ;
    wire \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_13 ;
    wire \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_14 ;
    wire \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_15 ;
    wire \current_shift_inst.un4_control_input_cry_16 ;
    wire \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ;
    wire bfn_11_18_0_;
    wire \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_17 ;
    wire \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_18 ;
    wire \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_19 ;
    wire \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ;
    wire \current_shift_inst.un4_control_input_cry_20 ;
    wire \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ;
    wire \current_shift_inst.un4_control_input_cry_21 ;
    wire \current_shift_inst.un4_control_input_cry_22 ;
    wire \current_shift_inst.un4_control_input_cry_23 ;
    wire \current_shift_inst.un4_control_input_cry_24 ;
    wire bfn_11_19_0_;
    wire \current_shift_inst.un4_control_input_cry_25 ;
    wire \current_shift_inst.un4_control_input_cry_26 ;
    wire \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ;
    wire \current_shift_inst.un4_control_input_cry_27 ;
    wire \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ;
    wire \current_shift_inst.un4_control_input_cry_28 ;
    wire \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ;
    wire \current_shift_inst.un4_control_input_cry_29 ;
    wire \current_shift_inst.un4_control_input_cry_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ;
    wire \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ;
    wire \current_shift_inst.z_31 ;
    wire \current_shift_inst.z_i_31 ;
    wire \current_shift_inst.elapsed_time_ns_phase_24 ;
    wire \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_phase_30 ;
    wire \current_shift_inst.elapsed_time_ns_phase_31 ;
    wire \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ;
    wire \current_shift_inst.un38_control_input_0_axb_31 ;
    wire \current_shift_inst.elapsed_time_ns_phase_26 ;
    wire \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ;
    wire \current_shift_inst.elapsed_time_ns_phase_22 ;
    wire \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ;
    wire \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ;
    wire il_max_comp1_D1;
    wire \phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_12_7_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire bfn_12_8_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire bfn_12_9_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ;
    wire \current_shift_inst.S3_sync_prevZ0 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt15 ;
    wire \current_shift_inst.S3_riseZ0 ;
    wire \current_shift_inst.S1_riseZ0 ;
    wire \current_shift_inst.N_199 ;
    wire \current_shift_inst.meas_stateZ0Z_0 ;
    wire measured_delay_hc_28;
    wire measured_delay_hc_29;
    wire measured_delay_hc_30;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ;
    wire bfn_12_14_0_;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_12_15_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_12_16_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_12_17_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.N_187_i_g ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input_axb_29 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input_axb_28 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input_axb_20 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input_axb_30 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input_axb_19 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input_axb_26 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input_axb_27 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input_axb_25 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un4_control_input_axb_22 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_12_19_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_12_20_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_12_21_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_12_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_191_i ;
    wire \current_shift_inst.timer_phase.N_188_i ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire il_max_comp2_c;
    wire il_max_comp2_D1;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire measured_delay_hc_25;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire measured_delay_hc_26;
    wire measured_delay_hc_24;
    wire s1_phy_c;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \delay_measurement_inst.prev_hc_sigZ0 ;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.N_221_0 ;
    wire \current_shift_inst.S3_syncZ0Z1 ;
    wire \current_shift_inst.S3_syncZ0Z0 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input_axb_24 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input_axb_15 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input_axb_16 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input_axb_17 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un4_control_input_axb_21 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.un4_control_input_axb_10 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un4_control_input_axb_11 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input_axb_12 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un4_control_input_axb_18 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input_axb_13 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un4_control_input_axb_14 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input_axb_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_321_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3 ;
    wire \delay_measurement_inst.delay_tr_timer.N_320_4 ;
    wire \delay_measurement_inst.N_305_1_cascade_ ;
    wire \delay_measurement_inst.N_305_1 ;
    wire \delay_measurement_inst.delay_tr_timer.N_299 ;
    wire \delay_measurement_inst.N_358_cascade_ ;
    wire \current_shift_inst.stop_timer_phaseZ0 ;
    wire \current_shift_inst.start_timer_phaseZ0 ;
    wire \current_shift_inst.timer_phase.runningZ0 ;
    wire \current_shift_inst.timer_phase.N_192_i ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ;
    wire \delay_measurement_inst.delay_tr_timer.N_296 ;
    wire \delay_measurement_inst.delay_tr_timer.N_293_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ;
    wire \delay_measurement_inst.N_307 ;
    wire s2_phy_c;
    wire \delay_measurement_inst.delay_hc_timer.N_335_i ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_14_5_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire bfn_14_6_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire bfn_14_7_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_N_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1 ;
    wire delay_hc_d2;
    wire \phase_controller_inst1.stoper_hc.time_passed11 ;
    wire \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.stateZ0Z_3 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire measured_delay_hc_18;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_2 ;
    wire red_c_i;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.N_232 ;
    wire \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_slave.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_slave.N_214 ;
    wire s4_phy_c;
    wire \phase_controller_slave.stateZ0Z_2 ;
    wire \phase_controller_slave.hc_time_passed ;
    wire s3_phy_c;
    wire \phase_controller_slave.N_211_cascade_ ;
    wire \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_ ;
    wire \phase_controller_slave.tr_time_passed ;
    wire \phase_controller_slave.stateZ0Z_0 ;
    wire il_max_comp2_D2;
    wire \phase_controller_slave.N_211 ;
    wire \phase_controller_slave.stateZ0Z_3 ;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire \delay_measurement_inst.prev_tr_sigZ0 ;
    wire start_stop_c;
    wire shift_flag_start;
    wire \phase_controller_slave.stateZ0Z_4 ;
    wire \phase_controller_slave.N_213 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_ ;
    wire \phase_controller_slave.stateZ0Z_1 ;
    wire il_min_comp2_D2;
    wire \phase_controller_slave.start_timer_tr_0_sqmuxa ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6_cascade_ ;
    wire \delay_measurement_inst.N_358 ;
    wire \delay_measurement_inst.delay_tr_timer.N_331 ;
    wire \delay_measurement_inst.delay_tr_timer.N_331_cascade_ ;
    wire \delay_measurement_inst.N_333_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.N_333 ;
    wire \delay_measurement_inst.N_328 ;
    wire \delay_measurement_inst.N_324 ;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire bfn_14_20_0_;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_reg3lto6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_reg3lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire bfn_14_21_0_;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire bfn_14_22_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_14_23_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.N_337_i ;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire delay_tr_d2;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.N_228 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire measured_delay_hc_11;
    wire measured_delay_hc_12;
    wire measured_delay_hc_19;
    wire measured_delay_hc_17;
    wire measured_delay_hc_9;
    wire measured_delay_hc_0;
    wire measured_delay_hc_6;
    wire measured_delay_hc_1;
    wire measured_delay_hc_3;
    wire measured_delay_hc_4;
    wire measured_delay_hc_16;
    wire measured_delay_hc_14;
    wire measured_delay_hc_10;
    wire measured_delay_hc_8;
    wire measured_delay_hc_31;
    wire measured_delay_hc_5;
    wire \phase_controller_inst1.stoper_hc.un1_startlt31_0 ;
    wire measured_delay_hc_13;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire measured_delay_hc_7;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0 ;
    wire \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ;
    wire bfn_15_13_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_15_14_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_15_15_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire \delay_measurement_inst.delay_tr_reg3lto14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_15_19_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_15_20_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_15_21_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_15_22_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_338_i ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_5_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_reg3lt31_0 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_6 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_16_11_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_8 ;
    wire bfn_16_12_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_16 ;
    wire bfn_16_13_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire \phase_controller_slave.stoper_tr.time_passed11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \delay_measurement_inst.N_284_1 ;
    wire \delay_measurement_inst.delay_tr_reg3lto15 ;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire measured_delay_tr_8;
    wire measured_delay_tr_2;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ;
    wire measured_delay_tr_1;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_20_li ;
    wire measured_delay_tr_3;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_1 ;
    wire bfn_16_18_0_;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_9 ;
    wire bfn_16_19_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_17 ;
    wire bfn_16_20_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_19 ;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_reg3lto31_0_0 ;
    wire measured_delay_hc_2;
    wire \delay_measurement_inst.un1_elapsed_time_hc ;
    wire \delay_measurement_inst.delay_hc_reg3 ;
    wire measured_delay_hc_15;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire bfn_17_8_0_;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_reg3lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_reg3lto9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire bfn_17_9_0_;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_reg3lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_reg3lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.N_335_i_g ;
    wire \phase_controller_slave.start_timer_hcZ0 ;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \phase_controller_inst1.N_231 ;
    wire \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_ ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_17_15_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_17_16_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_17_17_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_4 ;
    wire measured_delay_tr_7;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_7 ;
    wire measured_delay_tr_14;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_16 ;
    wire measured_delay_tr_6;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_ ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_10 ;
    wire measured_delay_tr_11;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_11 ;
    wire measured_delay_tr_12;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_12 ;
    wire measured_delay_tr_13;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ;
    wire measured_delay_tr_15;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ;
    wire measured_delay_tr_10;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_18_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_18_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_18_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_18_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_336_i ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_18_11_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire bfn_18_12_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire bfn_18_13_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.stoper_hc.time_passed11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire bfn_18_14_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire bfn_18_15_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire bfn_18_16_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.start_timer_trZ0 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire clk_100mhz_0;
    wire red_c_g;
    wire measured_delay_tr_18;
    wire measured_delay_tr_17;
    wire measured_delay_tr_19;
    wire measured_delay_tr_16;
    wire measured_delay_tr_5;
    wire measured_delay_tr_4;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_21 ;
    wire measured_delay_tr_9;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2 ;
    wire _gnd_net_;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__32628),
            .RESETB(N__34797),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__27778),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__27709),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__18556,N__18560,N__18557,N__18561,N__18558,N__18605,N__18584,N__18260,N__20513,N__18242,N__18451,N__18349,N__18399,N__18417,N__18380}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__27715,N__27712,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__27710,N__27714,N__27711,N__27713}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__27834),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__27830),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64}),
            .ADDSUBBOT(),
            .A({dangling_wire_65,N__18533,N__18526,N__18531,N__18525,N__18532,N__18524,N__18534,N__18521,N__18527,N__18520,N__18528,N__18522,N__18529,N__18523,N__18530}),
            .C({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .B({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,N__27837,N__27833,dangling_wire_89,dangling_wire_90,dangling_wire_91,N__27831,N__27836,N__27832,N__27835}),
            .OHOLDTOP(),
            .O({dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__48094),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__48096),
            .DIN(N__48095),
            .DOUT(N__48094),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__48096),
            .PADOUT(N__48095),
            .PADIN(N__48094),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__48085),
            .DIN(N__48084),
            .DOUT(N__48083),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__48085),
            .PADOUT(N__48084),
            .PADIN(N__48083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__48076),
            .DIN(N__48075),
            .DOUT(N__48074),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__48076),
            .PADOUT(N__48075),
            .PADIN(N__48074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__48067),
            .DIN(N__48066),
            .DOUT(N__48065),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__48067),
            .PADOUT(N__48066),
            .PADIN(N__48065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23682),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__48058),
            .DIN(N__48057),
            .DOUT(N__48056),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__48058),
            .PADOUT(N__48057),
            .PADIN(N__48056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__48049),
            .DIN(N__48048),
            .DOUT(N__48047),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__48049),
            .PADOUT(N__48048),
            .PADIN(N__48047),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33861),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__48040),
            .DIN(N__48039),
            .DOUT(N__48038),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__48040),
            .PADOUT(N__48039),
            .PADIN(N__48038),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__48031),
            .DIN(N__48030),
            .DOUT(N__48029),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__48031),
            .PADOUT(N__48030),
            .PADIN(N__48029),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__48022),
            .DIN(N__48021),
            .DOUT(N__48020),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__48022),
            .PADOUT(N__48021),
            .PADIN(N__48020),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__48013),
            .DIN(N__48012),
            .DOUT(N__48011),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__48013),
            .PADOUT(N__48012),
            .PADIN(N__48011),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32934),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__48004),
            .DIN(N__48003),
            .DOUT(N__48002),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__48004),
            .PADOUT(N__48003),
            .PADIN(N__48002),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34902),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__47995),
            .DIN(N__47994),
            .DOUT(N__47993),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__47995),
            .PADOUT(N__47994),
            .PADIN(N__47993),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__47986),
            .DIN(N__47985),
            .DOUT(N__47984),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__47986),
            .PADOUT(N__47985),
            .PADIN(N__47984),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34836),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11450 (
            .O(N__47967),
            .I(N__47964));
    LocalMux I__11449 (
            .O(N__47964),
            .I(N__47961));
    Odrv4 I__11448 (
            .O(N__47961),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__11447 (
            .O(N__47958),
            .I(N__47954));
    InMux I__11446 (
            .O(N__47957),
            .I(N__47951));
    LocalMux I__11445 (
            .O(N__47954),
            .I(N__47948));
    LocalMux I__11444 (
            .O(N__47951),
            .I(N__47945));
    Odrv12 I__11443 (
            .O(N__47948),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__11442 (
            .O(N__47945),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__11441 (
            .O(N__47940),
            .I(N__47933));
    CascadeMux I__11440 (
            .O(N__47939),
            .I(N__47927));
    CascadeMux I__11439 (
            .O(N__47938),
            .I(N__47918));
    CascadeMux I__11438 (
            .O(N__47937),
            .I(N__47915));
    CascadeMux I__11437 (
            .O(N__47936),
            .I(N__47912));
    InMux I__11436 (
            .O(N__47933),
            .I(N__47901));
    InMux I__11435 (
            .O(N__47932),
            .I(N__47901));
    CascadeMux I__11434 (
            .O(N__47931),
            .I(N__47896));
    CascadeMux I__11433 (
            .O(N__47930),
            .I(N__47893));
    InMux I__11432 (
            .O(N__47927),
            .I(N__47886));
    InMux I__11431 (
            .O(N__47926),
            .I(N__47886));
    InMux I__11430 (
            .O(N__47925),
            .I(N__47883));
    InMux I__11429 (
            .O(N__47924),
            .I(N__47880));
    InMux I__11428 (
            .O(N__47923),
            .I(N__47867));
    InMux I__11427 (
            .O(N__47922),
            .I(N__47867));
    InMux I__11426 (
            .O(N__47921),
            .I(N__47867));
    InMux I__11425 (
            .O(N__47918),
            .I(N__47867));
    InMux I__11424 (
            .O(N__47915),
            .I(N__47867));
    InMux I__11423 (
            .O(N__47912),
            .I(N__47867));
    InMux I__11422 (
            .O(N__47911),
            .I(N__47854));
    InMux I__11421 (
            .O(N__47910),
            .I(N__47854));
    InMux I__11420 (
            .O(N__47909),
            .I(N__47854));
    InMux I__11419 (
            .O(N__47908),
            .I(N__47854));
    InMux I__11418 (
            .O(N__47907),
            .I(N__47854));
    InMux I__11417 (
            .O(N__47906),
            .I(N__47854));
    LocalMux I__11416 (
            .O(N__47901),
            .I(N__47851));
    InMux I__11415 (
            .O(N__47900),
            .I(N__47848));
    CascadeMux I__11414 (
            .O(N__47899),
            .I(N__47845));
    InMux I__11413 (
            .O(N__47896),
            .I(N__47836));
    InMux I__11412 (
            .O(N__47893),
            .I(N__47836));
    InMux I__11411 (
            .O(N__47892),
            .I(N__47836));
    InMux I__11410 (
            .O(N__47891),
            .I(N__47836));
    LocalMux I__11409 (
            .O(N__47886),
            .I(N__47833));
    LocalMux I__11408 (
            .O(N__47883),
            .I(N__47830));
    LocalMux I__11407 (
            .O(N__47880),
            .I(N__47823));
    LocalMux I__11406 (
            .O(N__47867),
            .I(N__47823));
    LocalMux I__11405 (
            .O(N__47854),
            .I(N__47823));
    Span4Mux_v I__11404 (
            .O(N__47851),
            .I(N__47820));
    LocalMux I__11403 (
            .O(N__47848),
            .I(N__47817));
    InMux I__11402 (
            .O(N__47845),
            .I(N__47814));
    LocalMux I__11401 (
            .O(N__47836),
            .I(N__47809));
    Span4Mux_v I__11400 (
            .O(N__47833),
            .I(N__47809));
    Span4Mux_v I__11399 (
            .O(N__47830),
            .I(N__47804));
    Span4Mux_v I__11398 (
            .O(N__47823),
            .I(N__47804));
    Span4Mux_h I__11397 (
            .O(N__47820),
            .I(N__47799));
    Span4Mux_h I__11396 (
            .O(N__47817),
            .I(N__47799));
    LocalMux I__11395 (
            .O(N__47814),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__11394 (
            .O(N__47809),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__11393 (
            .O(N__47804),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__11392 (
            .O(N__47799),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__11391 (
            .O(N__47790),
            .I(N__47786));
    InMux I__11390 (
            .O(N__47789),
            .I(N__47759));
    InMux I__11389 (
            .O(N__47786),
            .I(N__47759));
    InMux I__11388 (
            .O(N__47785),
            .I(N__47759));
    InMux I__11387 (
            .O(N__47784),
            .I(N__47759));
    InMux I__11386 (
            .O(N__47783),
            .I(N__47759));
    InMux I__11385 (
            .O(N__47782),
            .I(N__47759));
    InMux I__11384 (
            .O(N__47781),
            .I(N__47759));
    InMux I__11383 (
            .O(N__47780),
            .I(N__47744));
    InMux I__11382 (
            .O(N__47779),
            .I(N__47744));
    InMux I__11381 (
            .O(N__47778),
            .I(N__47744));
    InMux I__11380 (
            .O(N__47777),
            .I(N__47744));
    InMux I__11379 (
            .O(N__47776),
            .I(N__47744));
    InMux I__11378 (
            .O(N__47775),
            .I(N__47744));
    InMux I__11377 (
            .O(N__47774),
            .I(N__47744));
    LocalMux I__11376 (
            .O(N__47759),
            .I(N__47738));
    LocalMux I__11375 (
            .O(N__47744),
            .I(N__47735));
    CascadeMux I__11374 (
            .O(N__47743),
            .I(N__47731));
    InMux I__11373 (
            .O(N__47742),
            .I(N__47726));
    CascadeMux I__11372 (
            .O(N__47741),
            .I(N__47722));
    Span4Mux_h I__11371 (
            .O(N__47738),
            .I(N__47716));
    Span4Mux_v I__11370 (
            .O(N__47735),
            .I(N__47716));
    InMux I__11369 (
            .O(N__47734),
            .I(N__47713));
    InMux I__11368 (
            .O(N__47731),
            .I(N__47710));
    InMux I__11367 (
            .O(N__47730),
            .I(N__47705));
    InMux I__11366 (
            .O(N__47729),
            .I(N__47705));
    LocalMux I__11365 (
            .O(N__47726),
            .I(N__47702));
    InMux I__11364 (
            .O(N__47725),
            .I(N__47699));
    InMux I__11363 (
            .O(N__47722),
            .I(N__47696));
    InMux I__11362 (
            .O(N__47721),
            .I(N__47693));
    Span4Mux_v I__11361 (
            .O(N__47716),
            .I(N__47688));
    LocalMux I__11360 (
            .O(N__47713),
            .I(N__47688));
    LocalMux I__11359 (
            .O(N__47710),
            .I(N__47681));
    LocalMux I__11358 (
            .O(N__47705),
            .I(N__47681));
    Span4Mux_h I__11357 (
            .O(N__47702),
            .I(N__47676));
    LocalMux I__11356 (
            .O(N__47699),
            .I(N__47676));
    LocalMux I__11355 (
            .O(N__47696),
            .I(N__47669));
    LocalMux I__11354 (
            .O(N__47693),
            .I(N__47669));
    Span4Mux_h I__11353 (
            .O(N__47688),
            .I(N__47669));
    InMux I__11352 (
            .O(N__47687),
            .I(N__47664));
    InMux I__11351 (
            .O(N__47686),
            .I(N__47664));
    Span12Mux_h I__11350 (
            .O(N__47681),
            .I(N__47661));
    Span4Mux_v I__11349 (
            .O(N__47676),
            .I(N__47658));
    Span4Mux_v I__11348 (
            .O(N__47669),
            .I(N__47655));
    LocalMux I__11347 (
            .O(N__47664),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv12 I__11346 (
            .O(N__47661),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__11345 (
            .O(N__47658),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__11344 (
            .O(N__47655),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    CascadeMux I__11343 (
            .O(N__47646),
            .I(N__47643));
    InMux I__11342 (
            .O(N__47643),
            .I(N__47640));
    LocalMux I__11341 (
            .O(N__47640),
            .I(N__47637));
    Span4Mux_h I__11340 (
            .O(N__47637),
            .I(N__47634));
    Odrv4 I__11339 (
            .O(N__47634),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    CascadeMux I__11338 (
            .O(N__47631),
            .I(N__47617));
    CascadeMux I__11337 (
            .O(N__47630),
            .I(N__47612));
    CascadeMux I__11336 (
            .O(N__47629),
            .I(N__47609));
    CascadeMux I__11335 (
            .O(N__47628),
            .I(N__47606));
    InMux I__11334 (
            .O(N__47627),
            .I(N__47590));
    InMux I__11333 (
            .O(N__47626),
            .I(N__47590));
    InMux I__11332 (
            .O(N__47625),
            .I(N__47590));
    InMux I__11331 (
            .O(N__47624),
            .I(N__47590));
    InMux I__11330 (
            .O(N__47623),
            .I(N__47590));
    InMux I__11329 (
            .O(N__47622),
            .I(N__47590));
    InMux I__11328 (
            .O(N__47621),
            .I(N__47590));
    InMux I__11327 (
            .O(N__47620),
            .I(N__47585));
    InMux I__11326 (
            .O(N__47617),
            .I(N__47585));
    InMux I__11325 (
            .O(N__47616),
            .I(N__47574));
    InMux I__11324 (
            .O(N__47615),
            .I(N__47574));
    InMux I__11323 (
            .O(N__47612),
            .I(N__47574));
    InMux I__11322 (
            .O(N__47609),
            .I(N__47574));
    InMux I__11321 (
            .O(N__47606),
            .I(N__47574));
    InMux I__11320 (
            .O(N__47605),
            .I(N__47566));
    LocalMux I__11319 (
            .O(N__47590),
            .I(N__47563));
    LocalMux I__11318 (
            .O(N__47585),
            .I(N__47558));
    LocalMux I__11317 (
            .O(N__47574),
            .I(N__47558));
    InMux I__11316 (
            .O(N__47573),
            .I(N__47551));
    InMux I__11315 (
            .O(N__47572),
            .I(N__47551));
    InMux I__11314 (
            .O(N__47571),
            .I(N__47551));
    InMux I__11313 (
            .O(N__47570),
            .I(N__47546));
    InMux I__11312 (
            .O(N__47569),
            .I(N__47546));
    LocalMux I__11311 (
            .O(N__47566),
            .I(N__47543));
    Span4Mux_h I__11310 (
            .O(N__47563),
            .I(N__47537));
    Span4Mux_v I__11309 (
            .O(N__47558),
            .I(N__47537));
    LocalMux I__11308 (
            .O(N__47551),
            .I(N__47532));
    LocalMux I__11307 (
            .O(N__47546),
            .I(N__47527));
    Span4Mux_v I__11306 (
            .O(N__47543),
            .I(N__47527));
    InMux I__11305 (
            .O(N__47542),
            .I(N__47524));
    Span4Mux_v I__11304 (
            .O(N__47537),
            .I(N__47521));
    InMux I__11303 (
            .O(N__47536),
            .I(N__47518));
    CascadeMux I__11302 (
            .O(N__47535),
            .I(N__47515));
    Span4Mux_v I__11301 (
            .O(N__47532),
            .I(N__47511));
    Span4Mux_h I__11300 (
            .O(N__47527),
            .I(N__47506));
    LocalMux I__11299 (
            .O(N__47524),
            .I(N__47506));
    Sp12to4 I__11298 (
            .O(N__47521),
            .I(N__47501));
    LocalMux I__11297 (
            .O(N__47518),
            .I(N__47501));
    InMux I__11296 (
            .O(N__47515),
            .I(N__47496));
    InMux I__11295 (
            .O(N__47514),
            .I(N__47496));
    Span4Mux_h I__11294 (
            .O(N__47511),
            .I(N__47491));
    Span4Mux_v I__11293 (
            .O(N__47506),
            .I(N__47491));
    Span12Mux_h I__11292 (
            .O(N__47501),
            .I(N__47488));
    LocalMux I__11291 (
            .O(N__47496),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__11290 (
            .O(N__47491),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv12 I__11289 (
            .O(N__47488),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__11288 (
            .O(N__47481),
            .I(N__47477));
    InMux I__11287 (
            .O(N__47480),
            .I(N__47474));
    LocalMux I__11286 (
            .O(N__47477),
            .I(N__47471));
    LocalMux I__11285 (
            .O(N__47474),
            .I(N__47468));
    Odrv12 I__11284 (
            .O(N__47471),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__11283 (
            .O(N__47468),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    ClkMux I__11282 (
            .O(N__47463),
            .I(N__46992));
    ClkMux I__11281 (
            .O(N__47462),
            .I(N__46992));
    ClkMux I__11280 (
            .O(N__47461),
            .I(N__46992));
    ClkMux I__11279 (
            .O(N__47460),
            .I(N__46992));
    ClkMux I__11278 (
            .O(N__47459),
            .I(N__46992));
    ClkMux I__11277 (
            .O(N__47458),
            .I(N__46992));
    ClkMux I__11276 (
            .O(N__47457),
            .I(N__46992));
    ClkMux I__11275 (
            .O(N__47456),
            .I(N__46992));
    ClkMux I__11274 (
            .O(N__47455),
            .I(N__46992));
    ClkMux I__11273 (
            .O(N__47454),
            .I(N__46992));
    ClkMux I__11272 (
            .O(N__47453),
            .I(N__46992));
    ClkMux I__11271 (
            .O(N__47452),
            .I(N__46992));
    ClkMux I__11270 (
            .O(N__47451),
            .I(N__46992));
    ClkMux I__11269 (
            .O(N__47450),
            .I(N__46992));
    ClkMux I__11268 (
            .O(N__47449),
            .I(N__46992));
    ClkMux I__11267 (
            .O(N__47448),
            .I(N__46992));
    ClkMux I__11266 (
            .O(N__47447),
            .I(N__46992));
    ClkMux I__11265 (
            .O(N__47446),
            .I(N__46992));
    ClkMux I__11264 (
            .O(N__47445),
            .I(N__46992));
    ClkMux I__11263 (
            .O(N__47444),
            .I(N__46992));
    ClkMux I__11262 (
            .O(N__47443),
            .I(N__46992));
    ClkMux I__11261 (
            .O(N__47442),
            .I(N__46992));
    ClkMux I__11260 (
            .O(N__47441),
            .I(N__46992));
    ClkMux I__11259 (
            .O(N__47440),
            .I(N__46992));
    ClkMux I__11258 (
            .O(N__47439),
            .I(N__46992));
    ClkMux I__11257 (
            .O(N__47438),
            .I(N__46992));
    ClkMux I__11256 (
            .O(N__47437),
            .I(N__46992));
    ClkMux I__11255 (
            .O(N__47436),
            .I(N__46992));
    ClkMux I__11254 (
            .O(N__47435),
            .I(N__46992));
    ClkMux I__11253 (
            .O(N__47434),
            .I(N__46992));
    ClkMux I__11252 (
            .O(N__47433),
            .I(N__46992));
    ClkMux I__11251 (
            .O(N__47432),
            .I(N__46992));
    ClkMux I__11250 (
            .O(N__47431),
            .I(N__46992));
    ClkMux I__11249 (
            .O(N__47430),
            .I(N__46992));
    ClkMux I__11248 (
            .O(N__47429),
            .I(N__46992));
    ClkMux I__11247 (
            .O(N__47428),
            .I(N__46992));
    ClkMux I__11246 (
            .O(N__47427),
            .I(N__46992));
    ClkMux I__11245 (
            .O(N__47426),
            .I(N__46992));
    ClkMux I__11244 (
            .O(N__47425),
            .I(N__46992));
    ClkMux I__11243 (
            .O(N__47424),
            .I(N__46992));
    ClkMux I__11242 (
            .O(N__47423),
            .I(N__46992));
    ClkMux I__11241 (
            .O(N__47422),
            .I(N__46992));
    ClkMux I__11240 (
            .O(N__47421),
            .I(N__46992));
    ClkMux I__11239 (
            .O(N__47420),
            .I(N__46992));
    ClkMux I__11238 (
            .O(N__47419),
            .I(N__46992));
    ClkMux I__11237 (
            .O(N__47418),
            .I(N__46992));
    ClkMux I__11236 (
            .O(N__47417),
            .I(N__46992));
    ClkMux I__11235 (
            .O(N__47416),
            .I(N__46992));
    ClkMux I__11234 (
            .O(N__47415),
            .I(N__46992));
    ClkMux I__11233 (
            .O(N__47414),
            .I(N__46992));
    ClkMux I__11232 (
            .O(N__47413),
            .I(N__46992));
    ClkMux I__11231 (
            .O(N__47412),
            .I(N__46992));
    ClkMux I__11230 (
            .O(N__47411),
            .I(N__46992));
    ClkMux I__11229 (
            .O(N__47410),
            .I(N__46992));
    ClkMux I__11228 (
            .O(N__47409),
            .I(N__46992));
    ClkMux I__11227 (
            .O(N__47408),
            .I(N__46992));
    ClkMux I__11226 (
            .O(N__47407),
            .I(N__46992));
    ClkMux I__11225 (
            .O(N__47406),
            .I(N__46992));
    ClkMux I__11224 (
            .O(N__47405),
            .I(N__46992));
    ClkMux I__11223 (
            .O(N__47404),
            .I(N__46992));
    ClkMux I__11222 (
            .O(N__47403),
            .I(N__46992));
    ClkMux I__11221 (
            .O(N__47402),
            .I(N__46992));
    ClkMux I__11220 (
            .O(N__47401),
            .I(N__46992));
    ClkMux I__11219 (
            .O(N__47400),
            .I(N__46992));
    ClkMux I__11218 (
            .O(N__47399),
            .I(N__46992));
    ClkMux I__11217 (
            .O(N__47398),
            .I(N__46992));
    ClkMux I__11216 (
            .O(N__47397),
            .I(N__46992));
    ClkMux I__11215 (
            .O(N__47396),
            .I(N__46992));
    ClkMux I__11214 (
            .O(N__47395),
            .I(N__46992));
    ClkMux I__11213 (
            .O(N__47394),
            .I(N__46992));
    ClkMux I__11212 (
            .O(N__47393),
            .I(N__46992));
    ClkMux I__11211 (
            .O(N__47392),
            .I(N__46992));
    ClkMux I__11210 (
            .O(N__47391),
            .I(N__46992));
    ClkMux I__11209 (
            .O(N__47390),
            .I(N__46992));
    ClkMux I__11208 (
            .O(N__47389),
            .I(N__46992));
    ClkMux I__11207 (
            .O(N__47388),
            .I(N__46992));
    ClkMux I__11206 (
            .O(N__47387),
            .I(N__46992));
    ClkMux I__11205 (
            .O(N__47386),
            .I(N__46992));
    ClkMux I__11204 (
            .O(N__47385),
            .I(N__46992));
    ClkMux I__11203 (
            .O(N__47384),
            .I(N__46992));
    ClkMux I__11202 (
            .O(N__47383),
            .I(N__46992));
    ClkMux I__11201 (
            .O(N__47382),
            .I(N__46992));
    ClkMux I__11200 (
            .O(N__47381),
            .I(N__46992));
    ClkMux I__11199 (
            .O(N__47380),
            .I(N__46992));
    ClkMux I__11198 (
            .O(N__47379),
            .I(N__46992));
    ClkMux I__11197 (
            .O(N__47378),
            .I(N__46992));
    ClkMux I__11196 (
            .O(N__47377),
            .I(N__46992));
    ClkMux I__11195 (
            .O(N__47376),
            .I(N__46992));
    ClkMux I__11194 (
            .O(N__47375),
            .I(N__46992));
    ClkMux I__11193 (
            .O(N__47374),
            .I(N__46992));
    ClkMux I__11192 (
            .O(N__47373),
            .I(N__46992));
    ClkMux I__11191 (
            .O(N__47372),
            .I(N__46992));
    ClkMux I__11190 (
            .O(N__47371),
            .I(N__46992));
    ClkMux I__11189 (
            .O(N__47370),
            .I(N__46992));
    ClkMux I__11188 (
            .O(N__47369),
            .I(N__46992));
    ClkMux I__11187 (
            .O(N__47368),
            .I(N__46992));
    ClkMux I__11186 (
            .O(N__47367),
            .I(N__46992));
    ClkMux I__11185 (
            .O(N__47366),
            .I(N__46992));
    ClkMux I__11184 (
            .O(N__47365),
            .I(N__46992));
    ClkMux I__11183 (
            .O(N__47364),
            .I(N__46992));
    ClkMux I__11182 (
            .O(N__47363),
            .I(N__46992));
    ClkMux I__11181 (
            .O(N__47362),
            .I(N__46992));
    ClkMux I__11180 (
            .O(N__47361),
            .I(N__46992));
    ClkMux I__11179 (
            .O(N__47360),
            .I(N__46992));
    ClkMux I__11178 (
            .O(N__47359),
            .I(N__46992));
    ClkMux I__11177 (
            .O(N__47358),
            .I(N__46992));
    ClkMux I__11176 (
            .O(N__47357),
            .I(N__46992));
    ClkMux I__11175 (
            .O(N__47356),
            .I(N__46992));
    ClkMux I__11174 (
            .O(N__47355),
            .I(N__46992));
    ClkMux I__11173 (
            .O(N__47354),
            .I(N__46992));
    ClkMux I__11172 (
            .O(N__47353),
            .I(N__46992));
    ClkMux I__11171 (
            .O(N__47352),
            .I(N__46992));
    ClkMux I__11170 (
            .O(N__47351),
            .I(N__46992));
    ClkMux I__11169 (
            .O(N__47350),
            .I(N__46992));
    ClkMux I__11168 (
            .O(N__47349),
            .I(N__46992));
    ClkMux I__11167 (
            .O(N__47348),
            .I(N__46992));
    ClkMux I__11166 (
            .O(N__47347),
            .I(N__46992));
    ClkMux I__11165 (
            .O(N__47346),
            .I(N__46992));
    ClkMux I__11164 (
            .O(N__47345),
            .I(N__46992));
    ClkMux I__11163 (
            .O(N__47344),
            .I(N__46992));
    ClkMux I__11162 (
            .O(N__47343),
            .I(N__46992));
    ClkMux I__11161 (
            .O(N__47342),
            .I(N__46992));
    ClkMux I__11160 (
            .O(N__47341),
            .I(N__46992));
    ClkMux I__11159 (
            .O(N__47340),
            .I(N__46992));
    ClkMux I__11158 (
            .O(N__47339),
            .I(N__46992));
    ClkMux I__11157 (
            .O(N__47338),
            .I(N__46992));
    ClkMux I__11156 (
            .O(N__47337),
            .I(N__46992));
    ClkMux I__11155 (
            .O(N__47336),
            .I(N__46992));
    ClkMux I__11154 (
            .O(N__47335),
            .I(N__46992));
    ClkMux I__11153 (
            .O(N__47334),
            .I(N__46992));
    ClkMux I__11152 (
            .O(N__47333),
            .I(N__46992));
    ClkMux I__11151 (
            .O(N__47332),
            .I(N__46992));
    ClkMux I__11150 (
            .O(N__47331),
            .I(N__46992));
    ClkMux I__11149 (
            .O(N__47330),
            .I(N__46992));
    ClkMux I__11148 (
            .O(N__47329),
            .I(N__46992));
    ClkMux I__11147 (
            .O(N__47328),
            .I(N__46992));
    ClkMux I__11146 (
            .O(N__47327),
            .I(N__46992));
    ClkMux I__11145 (
            .O(N__47326),
            .I(N__46992));
    ClkMux I__11144 (
            .O(N__47325),
            .I(N__46992));
    ClkMux I__11143 (
            .O(N__47324),
            .I(N__46992));
    ClkMux I__11142 (
            .O(N__47323),
            .I(N__46992));
    ClkMux I__11141 (
            .O(N__47322),
            .I(N__46992));
    ClkMux I__11140 (
            .O(N__47321),
            .I(N__46992));
    ClkMux I__11139 (
            .O(N__47320),
            .I(N__46992));
    ClkMux I__11138 (
            .O(N__47319),
            .I(N__46992));
    ClkMux I__11137 (
            .O(N__47318),
            .I(N__46992));
    ClkMux I__11136 (
            .O(N__47317),
            .I(N__46992));
    ClkMux I__11135 (
            .O(N__47316),
            .I(N__46992));
    ClkMux I__11134 (
            .O(N__47315),
            .I(N__46992));
    ClkMux I__11133 (
            .O(N__47314),
            .I(N__46992));
    ClkMux I__11132 (
            .O(N__47313),
            .I(N__46992));
    ClkMux I__11131 (
            .O(N__47312),
            .I(N__46992));
    ClkMux I__11130 (
            .O(N__47311),
            .I(N__46992));
    ClkMux I__11129 (
            .O(N__47310),
            .I(N__46992));
    ClkMux I__11128 (
            .O(N__47309),
            .I(N__46992));
    ClkMux I__11127 (
            .O(N__47308),
            .I(N__46992));
    ClkMux I__11126 (
            .O(N__47307),
            .I(N__46992));
    GlobalMux I__11125 (
            .O(N__46992),
            .I(clk_100mhz_0));
    CascadeMux I__11124 (
            .O(N__46989),
            .I(N__46981));
    CascadeMux I__11123 (
            .O(N__46988),
            .I(N__46978));
    InMux I__11122 (
            .O(N__46987),
            .I(N__46974));
    InMux I__11121 (
            .O(N__46986),
            .I(N__46971));
    InMux I__11120 (
            .O(N__46985),
            .I(N__46968));
    InMux I__11119 (
            .O(N__46984),
            .I(N__46965));
    InMux I__11118 (
            .O(N__46981),
            .I(N__46962));
    InMux I__11117 (
            .O(N__46978),
            .I(N__46959));
    InMux I__11116 (
            .O(N__46977),
            .I(N__46956));
    LocalMux I__11115 (
            .O(N__46974),
            .I(N__46953));
    LocalMux I__11114 (
            .O(N__46971),
            .I(N__46950));
    LocalMux I__11113 (
            .O(N__46968),
            .I(N__46947));
    LocalMux I__11112 (
            .O(N__46965),
            .I(N__46897));
    LocalMux I__11111 (
            .O(N__46962),
            .I(N__46878));
    LocalMux I__11110 (
            .O(N__46959),
            .I(N__46869));
    LocalMux I__11109 (
            .O(N__46956),
            .I(N__46837));
    Glb2LocalMux I__11108 (
            .O(N__46953),
            .I(N__46521));
    Glb2LocalMux I__11107 (
            .O(N__46950),
            .I(N__46521));
    Glb2LocalMux I__11106 (
            .O(N__46947),
            .I(N__46521));
    SRMux I__11105 (
            .O(N__46946),
            .I(N__46521));
    SRMux I__11104 (
            .O(N__46945),
            .I(N__46521));
    SRMux I__11103 (
            .O(N__46944),
            .I(N__46521));
    SRMux I__11102 (
            .O(N__46943),
            .I(N__46521));
    SRMux I__11101 (
            .O(N__46942),
            .I(N__46521));
    SRMux I__11100 (
            .O(N__46941),
            .I(N__46521));
    SRMux I__11099 (
            .O(N__46940),
            .I(N__46521));
    SRMux I__11098 (
            .O(N__46939),
            .I(N__46521));
    SRMux I__11097 (
            .O(N__46938),
            .I(N__46521));
    SRMux I__11096 (
            .O(N__46937),
            .I(N__46521));
    SRMux I__11095 (
            .O(N__46936),
            .I(N__46521));
    SRMux I__11094 (
            .O(N__46935),
            .I(N__46521));
    SRMux I__11093 (
            .O(N__46934),
            .I(N__46521));
    SRMux I__11092 (
            .O(N__46933),
            .I(N__46521));
    SRMux I__11091 (
            .O(N__46932),
            .I(N__46521));
    SRMux I__11090 (
            .O(N__46931),
            .I(N__46521));
    SRMux I__11089 (
            .O(N__46930),
            .I(N__46521));
    SRMux I__11088 (
            .O(N__46929),
            .I(N__46521));
    SRMux I__11087 (
            .O(N__46928),
            .I(N__46521));
    SRMux I__11086 (
            .O(N__46927),
            .I(N__46521));
    SRMux I__11085 (
            .O(N__46926),
            .I(N__46521));
    SRMux I__11084 (
            .O(N__46925),
            .I(N__46521));
    SRMux I__11083 (
            .O(N__46924),
            .I(N__46521));
    SRMux I__11082 (
            .O(N__46923),
            .I(N__46521));
    SRMux I__11081 (
            .O(N__46922),
            .I(N__46521));
    SRMux I__11080 (
            .O(N__46921),
            .I(N__46521));
    SRMux I__11079 (
            .O(N__46920),
            .I(N__46521));
    SRMux I__11078 (
            .O(N__46919),
            .I(N__46521));
    SRMux I__11077 (
            .O(N__46918),
            .I(N__46521));
    SRMux I__11076 (
            .O(N__46917),
            .I(N__46521));
    SRMux I__11075 (
            .O(N__46916),
            .I(N__46521));
    SRMux I__11074 (
            .O(N__46915),
            .I(N__46521));
    SRMux I__11073 (
            .O(N__46914),
            .I(N__46521));
    SRMux I__11072 (
            .O(N__46913),
            .I(N__46521));
    SRMux I__11071 (
            .O(N__46912),
            .I(N__46521));
    SRMux I__11070 (
            .O(N__46911),
            .I(N__46521));
    SRMux I__11069 (
            .O(N__46910),
            .I(N__46521));
    SRMux I__11068 (
            .O(N__46909),
            .I(N__46521));
    SRMux I__11067 (
            .O(N__46908),
            .I(N__46521));
    SRMux I__11066 (
            .O(N__46907),
            .I(N__46521));
    SRMux I__11065 (
            .O(N__46906),
            .I(N__46521));
    SRMux I__11064 (
            .O(N__46905),
            .I(N__46521));
    SRMux I__11063 (
            .O(N__46904),
            .I(N__46521));
    SRMux I__11062 (
            .O(N__46903),
            .I(N__46521));
    SRMux I__11061 (
            .O(N__46902),
            .I(N__46521));
    SRMux I__11060 (
            .O(N__46901),
            .I(N__46521));
    SRMux I__11059 (
            .O(N__46900),
            .I(N__46521));
    Glb2LocalMux I__11058 (
            .O(N__46897),
            .I(N__46521));
    SRMux I__11057 (
            .O(N__46896),
            .I(N__46521));
    SRMux I__11056 (
            .O(N__46895),
            .I(N__46521));
    SRMux I__11055 (
            .O(N__46894),
            .I(N__46521));
    SRMux I__11054 (
            .O(N__46893),
            .I(N__46521));
    SRMux I__11053 (
            .O(N__46892),
            .I(N__46521));
    SRMux I__11052 (
            .O(N__46891),
            .I(N__46521));
    SRMux I__11051 (
            .O(N__46890),
            .I(N__46521));
    SRMux I__11050 (
            .O(N__46889),
            .I(N__46521));
    SRMux I__11049 (
            .O(N__46888),
            .I(N__46521));
    SRMux I__11048 (
            .O(N__46887),
            .I(N__46521));
    SRMux I__11047 (
            .O(N__46886),
            .I(N__46521));
    SRMux I__11046 (
            .O(N__46885),
            .I(N__46521));
    SRMux I__11045 (
            .O(N__46884),
            .I(N__46521));
    SRMux I__11044 (
            .O(N__46883),
            .I(N__46521));
    SRMux I__11043 (
            .O(N__46882),
            .I(N__46521));
    SRMux I__11042 (
            .O(N__46881),
            .I(N__46521));
    Glb2LocalMux I__11041 (
            .O(N__46878),
            .I(N__46521));
    SRMux I__11040 (
            .O(N__46877),
            .I(N__46521));
    SRMux I__11039 (
            .O(N__46876),
            .I(N__46521));
    SRMux I__11038 (
            .O(N__46875),
            .I(N__46521));
    SRMux I__11037 (
            .O(N__46874),
            .I(N__46521));
    SRMux I__11036 (
            .O(N__46873),
            .I(N__46521));
    SRMux I__11035 (
            .O(N__46872),
            .I(N__46521));
    Glb2LocalMux I__11034 (
            .O(N__46869),
            .I(N__46521));
    SRMux I__11033 (
            .O(N__46868),
            .I(N__46521));
    SRMux I__11032 (
            .O(N__46867),
            .I(N__46521));
    SRMux I__11031 (
            .O(N__46866),
            .I(N__46521));
    SRMux I__11030 (
            .O(N__46865),
            .I(N__46521));
    SRMux I__11029 (
            .O(N__46864),
            .I(N__46521));
    SRMux I__11028 (
            .O(N__46863),
            .I(N__46521));
    SRMux I__11027 (
            .O(N__46862),
            .I(N__46521));
    SRMux I__11026 (
            .O(N__46861),
            .I(N__46521));
    SRMux I__11025 (
            .O(N__46860),
            .I(N__46521));
    SRMux I__11024 (
            .O(N__46859),
            .I(N__46521));
    SRMux I__11023 (
            .O(N__46858),
            .I(N__46521));
    SRMux I__11022 (
            .O(N__46857),
            .I(N__46521));
    SRMux I__11021 (
            .O(N__46856),
            .I(N__46521));
    SRMux I__11020 (
            .O(N__46855),
            .I(N__46521));
    SRMux I__11019 (
            .O(N__46854),
            .I(N__46521));
    SRMux I__11018 (
            .O(N__46853),
            .I(N__46521));
    SRMux I__11017 (
            .O(N__46852),
            .I(N__46521));
    SRMux I__11016 (
            .O(N__46851),
            .I(N__46521));
    SRMux I__11015 (
            .O(N__46850),
            .I(N__46521));
    SRMux I__11014 (
            .O(N__46849),
            .I(N__46521));
    SRMux I__11013 (
            .O(N__46848),
            .I(N__46521));
    SRMux I__11012 (
            .O(N__46847),
            .I(N__46521));
    SRMux I__11011 (
            .O(N__46846),
            .I(N__46521));
    SRMux I__11010 (
            .O(N__46845),
            .I(N__46521));
    SRMux I__11009 (
            .O(N__46844),
            .I(N__46521));
    SRMux I__11008 (
            .O(N__46843),
            .I(N__46521));
    SRMux I__11007 (
            .O(N__46842),
            .I(N__46521));
    SRMux I__11006 (
            .O(N__46841),
            .I(N__46521));
    SRMux I__11005 (
            .O(N__46840),
            .I(N__46521));
    Glb2LocalMux I__11004 (
            .O(N__46837),
            .I(N__46521));
    SRMux I__11003 (
            .O(N__46836),
            .I(N__46521));
    SRMux I__11002 (
            .O(N__46835),
            .I(N__46521));
    SRMux I__11001 (
            .O(N__46834),
            .I(N__46521));
    SRMux I__11000 (
            .O(N__46833),
            .I(N__46521));
    SRMux I__10999 (
            .O(N__46832),
            .I(N__46521));
    SRMux I__10998 (
            .O(N__46831),
            .I(N__46521));
    SRMux I__10997 (
            .O(N__46830),
            .I(N__46521));
    SRMux I__10996 (
            .O(N__46829),
            .I(N__46521));
    SRMux I__10995 (
            .O(N__46828),
            .I(N__46521));
    SRMux I__10994 (
            .O(N__46827),
            .I(N__46521));
    SRMux I__10993 (
            .O(N__46826),
            .I(N__46521));
    SRMux I__10992 (
            .O(N__46825),
            .I(N__46521));
    SRMux I__10991 (
            .O(N__46824),
            .I(N__46521));
    SRMux I__10990 (
            .O(N__46823),
            .I(N__46521));
    SRMux I__10989 (
            .O(N__46822),
            .I(N__46521));
    SRMux I__10988 (
            .O(N__46821),
            .I(N__46521));
    SRMux I__10987 (
            .O(N__46820),
            .I(N__46521));
    SRMux I__10986 (
            .O(N__46819),
            .I(N__46521));
    SRMux I__10985 (
            .O(N__46818),
            .I(N__46521));
    SRMux I__10984 (
            .O(N__46817),
            .I(N__46521));
    SRMux I__10983 (
            .O(N__46816),
            .I(N__46521));
    SRMux I__10982 (
            .O(N__46815),
            .I(N__46521));
    SRMux I__10981 (
            .O(N__46814),
            .I(N__46521));
    SRMux I__10980 (
            .O(N__46813),
            .I(N__46521));
    SRMux I__10979 (
            .O(N__46812),
            .I(N__46521));
    SRMux I__10978 (
            .O(N__46811),
            .I(N__46521));
    SRMux I__10977 (
            .O(N__46810),
            .I(N__46521));
    SRMux I__10976 (
            .O(N__46809),
            .I(N__46521));
    SRMux I__10975 (
            .O(N__46808),
            .I(N__46521));
    SRMux I__10974 (
            .O(N__46807),
            .I(N__46521));
    SRMux I__10973 (
            .O(N__46806),
            .I(N__46521));
    SRMux I__10972 (
            .O(N__46805),
            .I(N__46521));
    SRMux I__10971 (
            .O(N__46804),
            .I(N__46521));
    SRMux I__10970 (
            .O(N__46803),
            .I(N__46521));
    SRMux I__10969 (
            .O(N__46802),
            .I(N__46521));
    GlobalMux I__10968 (
            .O(N__46521),
            .I(N__46518));
    gio2CtrlBuf I__10967 (
            .O(N__46518),
            .I(red_c_g));
    InMux I__10966 (
            .O(N__46515),
            .I(N__46511));
    InMux I__10965 (
            .O(N__46514),
            .I(N__46507));
    LocalMux I__10964 (
            .O(N__46511),
            .I(N__46503));
    InMux I__10963 (
            .O(N__46510),
            .I(N__46500));
    LocalMux I__10962 (
            .O(N__46507),
            .I(N__46497));
    InMux I__10961 (
            .O(N__46506),
            .I(N__46494));
    Span4Mux_v I__10960 (
            .O(N__46503),
            .I(N__46489));
    LocalMux I__10959 (
            .O(N__46500),
            .I(N__46489));
    Span4Mux_h I__10958 (
            .O(N__46497),
            .I(N__46484));
    LocalMux I__10957 (
            .O(N__46494),
            .I(N__46484));
    Span4Mux_h I__10956 (
            .O(N__46489),
            .I(N__46481));
    Span4Mux_h I__10955 (
            .O(N__46484),
            .I(N__46478));
    Odrv4 I__10954 (
            .O(N__46481),
            .I(measured_delay_tr_18));
    Odrv4 I__10953 (
            .O(N__46478),
            .I(measured_delay_tr_18));
    InMux I__10952 (
            .O(N__46473),
            .I(N__46467));
    InMux I__10951 (
            .O(N__46472),
            .I(N__46464));
    InMux I__10950 (
            .O(N__46471),
            .I(N__46461));
    InMux I__10949 (
            .O(N__46470),
            .I(N__46458));
    LocalMux I__10948 (
            .O(N__46467),
            .I(N__46455));
    LocalMux I__10947 (
            .O(N__46464),
            .I(N__46452));
    LocalMux I__10946 (
            .O(N__46461),
            .I(N__46447));
    LocalMux I__10945 (
            .O(N__46458),
            .I(N__46447));
    Span4Mux_v I__10944 (
            .O(N__46455),
            .I(N__46440));
    Span4Mux_v I__10943 (
            .O(N__46452),
            .I(N__46440));
    Span4Mux_h I__10942 (
            .O(N__46447),
            .I(N__46440));
    Span4Mux_h I__10941 (
            .O(N__46440),
            .I(N__46437));
    Odrv4 I__10940 (
            .O(N__46437),
            .I(measured_delay_tr_17));
    CascadeMux I__10939 (
            .O(N__46434),
            .I(N__46429));
    InMux I__10938 (
            .O(N__46433),
            .I(N__46426));
    CascadeMux I__10937 (
            .O(N__46432),
            .I(N__46423));
    InMux I__10936 (
            .O(N__46429),
            .I(N__46419));
    LocalMux I__10935 (
            .O(N__46426),
            .I(N__46416));
    InMux I__10934 (
            .O(N__46423),
            .I(N__46413));
    InMux I__10933 (
            .O(N__46422),
            .I(N__46410));
    LocalMux I__10932 (
            .O(N__46419),
            .I(N__46407));
    Span4Mux_v I__10931 (
            .O(N__46416),
            .I(N__46402));
    LocalMux I__10930 (
            .O(N__46413),
            .I(N__46402));
    LocalMux I__10929 (
            .O(N__46410),
            .I(N__46397));
    Span4Mux_v I__10928 (
            .O(N__46407),
            .I(N__46397));
    Span4Mux_v I__10927 (
            .O(N__46402),
            .I(N__46394));
    Span4Mux_h I__10926 (
            .O(N__46397),
            .I(N__46391));
    Span4Mux_h I__10925 (
            .O(N__46394),
            .I(N__46388));
    Odrv4 I__10924 (
            .O(N__46391),
            .I(measured_delay_tr_19));
    Odrv4 I__10923 (
            .O(N__46388),
            .I(measured_delay_tr_19));
    InMux I__10922 (
            .O(N__46383),
            .I(N__46377));
    InMux I__10921 (
            .O(N__46382),
            .I(N__46374));
    InMux I__10920 (
            .O(N__46381),
            .I(N__46371));
    InMux I__10919 (
            .O(N__46380),
            .I(N__46368));
    LocalMux I__10918 (
            .O(N__46377),
            .I(N__46365));
    LocalMux I__10917 (
            .O(N__46374),
            .I(N__46362));
    LocalMux I__10916 (
            .O(N__46371),
            .I(N__46357));
    LocalMux I__10915 (
            .O(N__46368),
            .I(N__46357));
    Span4Mux_v I__10914 (
            .O(N__46365),
            .I(N__46350));
    Span4Mux_v I__10913 (
            .O(N__46362),
            .I(N__46350));
    Span4Mux_h I__10912 (
            .O(N__46357),
            .I(N__46350));
    Span4Mux_h I__10911 (
            .O(N__46350),
            .I(N__46347));
    Odrv4 I__10910 (
            .O(N__46347),
            .I(measured_delay_tr_16));
    CascadeMux I__10909 (
            .O(N__46344),
            .I(N__46341));
    InMux I__10908 (
            .O(N__46341),
            .I(N__46337));
    InMux I__10907 (
            .O(N__46340),
            .I(N__46333));
    LocalMux I__10906 (
            .O(N__46337),
            .I(N__46330));
    CascadeMux I__10905 (
            .O(N__46336),
            .I(N__46327));
    LocalMux I__10904 (
            .O(N__46333),
            .I(N__46324));
    Span4Mux_h I__10903 (
            .O(N__46330),
            .I(N__46321));
    InMux I__10902 (
            .O(N__46327),
            .I(N__46318));
    Span4Mux_v I__10901 (
            .O(N__46324),
            .I(N__46315));
    Odrv4 I__10900 (
            .O(N__46321),
            .I(measured_delay_tr_5));
    LocalMux I__10899 (
            .O(N__46318),
            .I(measured_delay_tr_5));
    Odrv4 I__10898 (
            .O(N__46315),
            .I(measured_delay_tr_5));
    InMux I__10897 (
            .O(N__46308),
            .I(N__46303));
    CascadeMux I__10896 (
            .O(N__46307),
            .I(N__46300));
    InMux I__10895 (
            .O(N__46306),
            .I(N__46297));
    LocalMux I__10894 (
            .O(N__46303),
            .I(N__46294));
    InMux I__10893 (
            .O(N__46300),
            .I(N__46291));
    LocalMux I__10892 (
            .O(N__46297),
            .I(N__46288));
    Span4Mux_h I__10891 (
            .O(N__46294),
            .I(N__46285));
    LocalMux I__10890 (
            .O(N__46291),
            .I(N__46280));
    Span4Mux_v I__10889 (
            .O(N__46288),
            .I(N__46280));
    Odrv4 I__10888 (
            .O(N__46285),
            .I(measured_delay_tr_4));
    Odrv4 I__10887 (
            .O(N__46280),
            .I(measured_delay_tr_4));
    CascadeMux I__10886 (
            .O(N__46275),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_ ));
    InMux I__10885 (
            .O(N__46272),
            .I(N__46268));
    InMux I__10884 (
            .O(N__46271),
            .I(N__46265));
    LocalMux I__10883 (
            .O(N__46268),
            .I(\phase_controller_inst1.stoper_tr.N_21 ));
    LocalMux I__10882 (
            .O(N__46265),
            .I(\phase_controller_inst1.stoper_tr.N_21 ));
    CascadeMux I__10881 (
            .O(N__46260),
            .I(N__46257));
    InMux I__10880 (
            .O(N__46257),
            .I(N__46252));
    InMux I__10879 (
            .O(N__46256),
            .I(N__46249));
    InMux I__10878 (
            .O(N__46255),
            .I(N__46245));
    LocalMux I__10877 (
            .O(N__46252),
            .I(N__46242));
    LocalMux I__10876 (
            .O(N__46249),
            .I(N__46239));
    InMux I__10875 (
            .O(N__46248),
            .I(N__46236));
    LocalMux I__10874 (
            .O(N__46245),
            .I(N__46233));
    Span4Mux_h I__10873 (
            .O(N__46242),
            .I(N__46230));
    Sp12to4 I__10872 (
            .O(N__46239),
            .I(N__46225));
    LocalMux I__10871 (
            .O(N__46236),
            .I(N__46225));
    Span4Mux_v I__10870 (
            .O(N__46233),
            .I(N__46222));
    Odrv4 I__10869 (
            .O(N__46230),
            .I(measured_delay_tr_9));
    Odrv12 I__10868 (
            .O(N__46225),
            .I(measured_delay_tr_9));
    Odrv4 I__10867 (
            .O(N__46222),
            .I(measured_delay_tr_9));
    InMux I__10866 (
            .O(N__46215),
            .I(N__46211));
    InMux I__10865 (
            .O(N__46214),
            .I(N__46208));
    LocalMux I__10864 (
            .O(N__46211),
            .I(N__46205));
    LocalMux I__10863 (
            .O(N__46208),
            .I(N__46202));
    Odrv12 I__10862 (
            .O(N__46205),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ));
    Odrv4 I__10861 (
            .O(N__46202),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ));
    CascadeMux I__10860 (
            .O(N__46197),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3_cascade_ ));
    InMux I__10859 (
            .O(N__46194),
            .I(N__46189));
    InMux I__10858 (
            .O(N__46193),
            .I(N__46186));
    InMux I__10857 (
            .O(N__46192),
            .I(N__46183));
    LocalMux I__10856 (
            .O(N__46189),
            .I(N__46180));
    LocalMux I__10855 (
            .O(N__46186),
            .I(N__46175));
    LocalMux I__10854 (
            .O(N__46183),
            .I(N__46175));
    Span4Mux_h I__10853 (
            .O(N__46180),
            .I(N__46171));
    Span4Mux_h I__10852 (
            .O(N__46175),
            .I(N__46168));
    InMux I__10851 (
            .O(N__46174),
            .I(N__46165));
    Odrv4 I__10850 (
            .O(N__46171),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ));
    Odrv4 I__10849 (
            .O(N__46168),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ));
    LocalMux I__10848 (
            .O(N__46165),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ));
    InMux I__10847 (
            .O(N__46158),
            .I(N__46148));
    InMux I__10846 (
            .O(N__46157),
            .I(N__46148));
    InMux I__10845 (
            .O(N__46156),
            .I(N__46148));
    InMux I__10844 (
            .O(N__46155),
            .I(N__46143));
    LocalMux I__10843 (
            .O(N__46148),
            .I(N__46140));
    InMux I__10842 (
            .O(N__46147),
            .I(N__46135));
    InMux I__10841 (
            .O(N__46146),
            .I(N__46135));
    LocalMux I__10840 (
            .O(N__46143),
            .I(N__46132));
    Span4Mux_v I__10839 (
            .O(N__46140),
            .I(N__46127));
    LocalMux I__10838 (
            .O(N__46135),
            .I(N__46127));
    Span4Mux_h I__10837 (
            .O(N__46132),
            .I(N__46124));
    Span4Mux_h I__10836 (
            .O(N__46127),
            .I(N__46121));
    Odrv4 I__10835 (
            .O(N__46124),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ));
    Odrv4 I__10834 (
            .O(N__46121),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ));
    InMux I__10833 (
            .O(N__46116),
            .I(N__46113));
    LocalMux I__10832 (
            .O(N__46113),
            .I(N__46110));
    Odrv4 I__10831 (
            .O(N__46110),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__10830 (
            .O(N__46107),
            .I(N__46104));
    LocalMux I__10829 (
            .O(N__46104),
            .I(N__46101));
    Odrv4 I__10828 (
            .O(N__46101),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__10827 (
            .O(N__46098),
            .I(N__46092));
    InMux I__10826 (
            .O(N__46097),
            .I(N__46092));
    LocalMux I__10825 (
            .O(N__46092),
            .I(N__46089));
    Odrv12 I__10824 (
            .O(N__46089),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2 ));
    CascadeMux I__10823 (
            .O(N__46086),
            .I(N__46083));
    InMux I__10822 (
            .O(N__46083),
            .I(N__46080));
    LocalMux I__10821 (
            .O(N__46080),
            .I(N__46077));
    Odrv12 I__10820 (
            .O(N__46077),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__10819 (
            .O(N__46074),
            .I(N__46071));
    LocalMux I__10818 (
            .O(N__46071),
            .I(N__46067));
    InMux I__10817 (
            .O(N__46070),
            .I(N__46064));
    Span4Mux_h I__10816 (
            .O(N__46067),
            .I(N__46059));
    LocalMux I__10815 (
            .O(N__46064),
            .I(N__46059));
    Odrv4 I__10814 (
            .O(N__46059),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__10813 (
            .O(N__46056),
            .I(N__46053));
    LocalMux I__10812 (
            .O(N__46053),
            .I(N__46050));
    Span4Mux_h I__10811 (
            .O(N__46050),
            .I(N__46047));
    Odrv4 I__10810 (
            .O(N__46047),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__10809 (
            .O(N__46044),
            .I(N__46040));
    InMux I__10808 (
            .O(N__46043),
            .I(N__46037));
    LocalMux I__10807 (
            .O(N__46040),
            .I(N__46034));
    LocalMux I__10806 (
            .O(N__46037),
            .I(N__46031));
    Odrv12 I__10805 (
            .O(N__46034),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__10804 (
            .O(N__46031),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__10803 (
            .O(N__46026),
            .I(N__46023));
    LocalMux I__10802 (
            .O(N__46023),
            .I(N__46020));
    Span4Mux_v I__10801 (
            .O(N__46020),
            .I(N__46017));
    Odrv4 I__10800 (
            .O(N__46017),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__10799 (
            .O(N__46014),
            .I(N__46010));
    InMux I__10798 (
            .O(N__46013),
            .I(N__46007));
    LocalMux I__10797 (
            .O(N__46010),
            .I(N__46002));
    LocalMux I__10796 (
            .O(N__46007),
            .I(N__46002));
    Odrv4 I__10795 (
            .O(N__46002),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__10794 (
            .O(N__45999),
            .I(N__45996));
    LocalMux I__10793 (
            .O(N__45996),
            .I(N__45991));
    InMux I__10792 (
            .O(N__45995),
            .I(N__45988));
    InMux I__10791 (
            .O(N__45994),
            .I(N__45984));
    Span4Mux_v I__10790 (
            .O(N__45991),
            .I(N__45979));
    LocalMux I__10789 (
            .O(N__45988),
            .I(N__45979));
    InMux I__10788 (
            .O(N__45987),
            .I(N__45976));
    LocalMux I__10787 (
            .O(N__45984),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    Odrv4 I__10786 (
            .O(N__45979),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    LocalMux I__10785 (
            .O(N__45976),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    InMux I__10784 (
            .O(N__45969),
            .I(N__45963));
    InMux I__10783 (
            .O(N__45968),
            .I(N__45963));
    LocalMux I__10782 (
            .O(N__45963),
            .I(N__45960));
    Span4Mux_h I__10781 (
            .O(N__45960),
            .I(N__45953));
    InMux I__10780 (
            .O(N__45959),
            .I(N__45948));
    InMux I__10779 (
            .O(N__45958),
            .I(N__45948));
    InMux I__10778 (
            .O(N__45957),
            .I(N__45945));
    InMux I__10777 (
            .O(N__45956),
            .I(N__45942));
    Span4Mux_v I__10776 (
            .O(N__45953),
            .I(N__45937));
    LocalMux I__10775 (
            .O(N__45948),
            .I(N__45937));
    LocalMux I__10774 (
            .O(N__45945),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__10773 (
            .O(N__45942),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__10772 (
            .O(N__45937),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__10771 (
            .O(N__45930),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    CascadeMux I__10770 (
            .O(N__45927),
            .I(N__45924));
    InMux I__10769 (
            .O(N__45924),
            .I(N__45919));
    InMux I__10768 (
            .O(N__45923),
            .I(N__45916));
    InMux I__10767 (
            .O(N__45922),
            .I(N__45913));
    LocalMux I__10766 (
            .O(N__45919),
            .I(N__45910));
    LocalMux I__10765 (
            .O(N__45916),
            .I(N__45907));
    LocalMux I__10764 (
            .O(N__45913),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__10763 (
            .O(N__45910),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__10762 (
            .O(N__45907),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__10761 (
            .O(N__45900),
            .I(N__45897));
    LocalMux I__10760 (
            .O(N__45897),
            .I(N__45894));
    Odrv4 I__10759 (
            .O(N__45894),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__10758 (
            .O(N__45891),
            .I(N__45887));
    InMux I__10757 (
            .O(N__45890),
            .I(N__45884));
    LocalMux I__10756 (
            .O(N__45887),
            .I(N__45881));
    LocalMux I__10755 (
            .O(N__45884),
            .I(N__45878));
    Odrv4 I__10754 (
            .O(N__45881),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__10753 (
            .O(N__45878),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__10752 (
            .O(N__45873),
            .I(N__45870));
    LocalMux I__10751 (
            .O(N__45870),
            .I(N__45867));
    Odrv4 I__10750 (
            .O(N__45867),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__10749 (
            .O(N__45864),
            .I(N__45860));
    InMux I__10748 (
            .O(N__45863),
            .I(N__45857));
    LocalMux I__10747 (
            .O(N__45860),
            .I(N__45854));
    LocalMux I__10746 (
            .O(N__45857),
            .I(N__45851));
    Odrv12 I__10745 (
            .O(N__45854),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__10744 (
            .O(N__45851),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__10743 (
            .O(N__45846),
            .I(N__45843));
    InMux I__10742 (
            .O(N__45843),
            .I(N__45840));
    LocalMux I__10741 (
            .O(N__45840),
            .I(N__45837));
    Odrv4 I__10740 (
            .O(N__45837),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__10739 (
            .O(N__45834),
            .I(N__45830));
    InMux I__10738 (
            .O(N__45833),
            .I(N__45827));
    LocalMux I__10737 (
            .O(N__45830),
            .I(N__45822));
    LocalMux I__10736 (
            .O(N__45827),
            .I(N__45822));
    Odrv4 I__10735 (
            .O(N__45822),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__10734 (
            .O(N__45819),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__10733 (
            .O(N__45816),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__10732 (
            .O(N__45813),
            .I(N__45810));
    LocalMux I__10731 (
            .O(N__45810),
            .I(N__45807));
    Odrv4 I__10730 (
            .O(N__45807),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ));
    CascadeMux I__10729 (
            .O(N__45804),
            .I(N__45801));
    InMux I__10728 (
            .O(N__45801),
            .I(N__45798));
    LocalMux I__10727 (
            .O(N__45798),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__10726 (
            .O(N__45795),
            .I(N__45791));
    InMux I__10725 (
            .O(N__45794),
            .I(N__45788));
    LocalMux I__10724 (
            .O(N__45791),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__10723 (
            .O(N__45788),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__10722 (
            .O(N__45783),
            .I(N__45780));
    LocalMux I__10721 (
            .O(N__45780),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    InMux I__10720 (
            .O(N__45777),
            .I(N__45773));
    InMux I__10719 (
            .O(N__45776),
            .I(N__45770));
    LocalMux I__10718 (
            .O(N__45773),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__10717 (
            .O(N__45770),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__10716 (
            .O(N__45765),
            .I(N__45762));
    LocalMux I__10715 (
            .O(N__45762),
            .I(N__45759));
    Span4Mux_v I__10714 (
            .O(N__45759),
            .I(N__45756));
    Odrv4 I__10713 (
            .O(N__45756),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ));
    CascadeMux I__10712 (
            .O(N__45753),
            .I(N__45745));
    CascadeMux I__10711 (
            .O(N__45752),
            .I(N__45742));
    CascadeMux I__10710 (
            .O(N__45751),
            .I(N__45735));
    CascadeMux I__10709 (
            .O(N__45750),
            .I(N__45727));
    CascadeMux I__10708 (
            .O(N__45749),
            .I(N__45720));
    CascadeMux I__10707 (
            .O(N__45748),
            .I(N__45717));
    InMux I__10706 (
            .O(N__45745),
            .I(N__45710));
    InMux I__10705 (
            .O(N__45742),
            .I(N__45710));
    InMux I__10704 (
            .O(N__45741),
            .I(N__45701));
    InMux I__10703 (
            .O(N__45740),
            .I(N__45701));
    InMux I__10702 (
            .O(N__45739),
            .I(N__45701));
    InMux I__10701 (
            .O(N__45738),
            .I(N__45701));
    InMux I__10700 (
            .O(N__45735),
            .I(N__45698));
    InMux I__10699 (
            .O(N__45734),
            .I(N__45691));
    InMux I__10698 (
            .O(N__45733),
            .I(N__45691));
    InMux I__10697 (
            .O(N__45732),
            .I(N__45691));
    InMux I__10696 (
            .O(N__45731),
            .I(N__45688));
    InMux I__10695 (
            .O(N__45730),
            .I(N__45685));
    InMux I__10694 (
            .O(N__45727),
            .I(N__45682));
    InMux I__10693 (
            .O(N__45726),
            .I(N__45675));
    InMux I__10692 (
            .O(N__45725),
            .I(N__45675));
    InMux I__10691 (
            .O(N__45724),
            .I(N__45675));
    InMux I__10690 (
            .O(N__45723),
            .I(N__45670));
    InMux I__10689 (
            .O(N__45720),
            .I(N__45661));
    InMux I__10688 (
            .O(N__45717),
            .I(N__45661));
    InMux I__10687 (
            .O(N__45716),
            .I(N__45661));
    InMux I__10686 (
            .O(N__45715),
            .I(N__45661));
    LocalMux I__10685 (
            .O(N__45710),
            .I(N__45651));
    LocalMux I__10684 (
            .O(N__45701),
            .I(N__45651));
    LocalMux I__10683 (
            .O(N__45698),
            .I(N__45651));
    LocalMux I__10682 (
            .O(N__45691),
            .I(N__45651));
    LocalMux I__10681 (
            .O(N__45688),
            .I(N__45648));
    LocalMux I__10680 (
            .O(N__45685),
            .I(N__45641));
    LocalMux I__10679 (
            .O(N__45682),
            .I(N__45641));
    LocalMux I__10678 (
            .O(N__45675),
            .I(N__45641));
    InMux I__10677 (
            .O(N__45674),
            .I(N__45636));
    InMux I__10676 (
            .O(N__45673),
            .I(N__45636));
    LocalMux I__10675 (
            .O(N__45670),
            .I(N__45633));
    LocalMux I__10674 (
            .O(N__45661),
            .I(N__45630));
    InMux I__10673 (
            .O(N__45660),
            .I(N__45627));
    Span4Mux_v I__10672 (
            .O(N__45651),
            .I(N__45624));
    Span12Mux_v I__10671 (
            .O(N__45648),
            .I(N__45621));
    Span12Mux_h I__10670 (
            .O(N__45641),
            .I(N__45618));
    LocalMux I__10669 (
            .O(N__45636),
            .I(N__45609));
    Span4Mux_v I__10668 (
            .O(N__45633),
            .I(N__45609));
    Span4Mux_h I__10667 (
            .O(N__45630),
            .I(N__45609));
    LocalMux I__10666 (
            .O(N__45627),
            .I(N__45609));
    Odrv4 I__10665 (
            .O(N__45624),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv12 I__10664 (
            .O(N__45621),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv12 I__10663 (
            .O(N__45618),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__10662 (
            .O(N__45609),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    CascadeMux I__10661 (
            .O(N__45600),
            .I(N__45593));
    CascadeMux I__10660 (
            .O(N__45599),
            .I(N__45587));
    CascadeMux I__10659 (
            .O(N__45598),
            .I(N__45584));
    CascadeMux I__10658 (
            .O(N__45597),
            .I(N__45580));
    CascadeMux I__10657 (
            .O(N__45596),
            .I(N__45577));
    InMux I__10656 (
            .O(N__45593),
            .I(N__45570));
    CascadeMux I__10655 (
            .O(N__45592),
            .I(N__45566));
    CascadeMux I__10654 (
            .O(N__45591),
            .I(N__45562));
    InMux I__10653 (
            .O(N__45590),
            .I(N__45553));
    InMux I__10652 (
            .O(N__45587),
            .I(N__45553));
    InMux I__10651 (
            .O(N__45584),
            .I(N__45544));
    InMux I__10650 (
            .O(N__45583),
            .I(N__45544));
    InMux I__10649 (
            .O(N__45580),
            .I(N__45544));
    InMux I__10648 (
            .O(N__45577),
            .I(N__45544));
    InMux I__10647 (
            .O(N__45576),
            .I(N__45535));
    InMux I__10646 (
            .O(N__45575),
            .I(N__45535));
    InMux I__10645 (
            .O(N__45574),
            .I(N__45535));
    InMux I__10644 (
            .O(N__45573),
            .I(N__45535));
    LocalMux I__10643 (
            .O(N__45570),
            .I(N__45530));
    InMux I__10642 (
            .O(N__45569),
            .I(N__45521));
    InMux I__10641 (
            .O(N__45566),
            .I(N__45521));
    InMux I__10640 (
            .O(N__45565),
            .I(N__45521));
    InMux I__10639 (
            .O(N__45562),
            .I(N__45521));
    CascadeMux I__10638 (
            .O(N__45561),
            .I(N__45518));
    CascadeMux I__10637 (
            .O(N__45560),
            .I(N__45514));
    CascadeMux I__10636 (
            .O(N__45559),
            .I(N__45510));
    CascadeMux I__10635 (
            .O(N__45558),
            .I(N__45507));
    LocalMux I__10634 (
            .O(N__45553),
            .I(N__45504));
    LocalMux I__10633 (
            .O(N__45544),
            .I(N__45499));
    LocalMux I__10632 (
            .O(N__45535),
            .I(N__45499));
    CascadeMux I__10631 (
            .O(N__45534),
            .I(N__45496));
    InMux I__10630 (
            .O(N__45533),
            .I(N__45492));
    Span4Mux_v I__10629 (
            .O(N__45530),
            .I(N__45489));
    LocalMux I__10628 (
            .O(N__45521),
            .I(N__45486));
    InMux I__10627 (
            .O(N__45518),
            .I(N__45473));
    InMux I__10626 (
            .O(N__45517),
            .I(N__45473));
    InMux I__10625 (
            .O(N__45514),
            .I(N__45473));
    InMux I__10624 (
            .O(N__45513),
            .I(N__45473));
    InMux I__10623 (
            .O(N__45510),
            .I(N__45473));
    InMux I__10622 (
            .O(N__45507),
            .I(N__45473));
    Span4Mux_v I__10621 (
            .O(N__45504),
            .I(N__45468));
    Span4Mux_v I__10620 (
            .O(N__45499),
            .I(N__45468));
    InMux I__10619 (
            .O(N__45496),
            .I(N__45463));
    InMux I__10618 (
            .O(N__45495),
            .I(N__45463));
    LocalMux I__10617 (
            .O(N__45492),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__10616 (
            .O(N__45489),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__10615 (
            .O(N__45486),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    LocalMux I__10614 (
            .O(N__45473),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__10613 (
            .O(N__45468),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    LocalMux I__10612 (
            .O(N__45463),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    InMux I__10611 (
            .O(N__45450),
            .I(N__45438));
    InMux I__10610 (
            .O(N__45449),
            .I(N__45429));
    InMux I__10609 (
            .O(N__45448),
            .I(N__45429));
    InMux I__10608 (
            .O(N__45447),
            .I(N__45429));
    InMux I__10607 (
            .O(N__45446),
            .I(N__45429));
    InMux I__10606 (
            .O(N__45445),
            .I(N__45420));
    InMux I__10605 (
            .O(N__45444),
            .I(N__45420));
    InMux I__10604 (
            .O(N__45443),
            .I(N__45420));
    InMux I__10603 (
            .O(N__45442),
            .I(N__45420));
    CascadeMux I__10602 (
            .O(N__45441),
            .I(N__45408));
    LocalMux I__10601 (
            .O(N__45438),
            .I(N__45402));
    LocalMux I__10600 (
            .O(N__45429),
            .I(N__45399));
    LocalMux I__10599 (
            .O(N__45420),
            .I(N__45396));
    InMux I__10598 (
            .O(N__45419),
            .I(N__45383));
    InMux I__10597 (
            .O(N__45418),
            .I(N__45383));
    InMux I__10596 (
            .O(N__45417),
            .I(N__45383));
    InMux I__10595 (
            .O(N__45416),
            .I(N__45383));
    InMux I__10594 (
            .O(N__45415),
            .I(N__45383));
    InMux I__10593 (
            .O(N__45414),
            .I(N__45383));
    CascadeMux I__10592 (
            .O(N__45413),
            .I(N__45380));
    InMux I__10591 (
            .O(N__45412),
            .I(N__45374));
    InMux I__10590 (
            .O(N__45411),
            .I(N__45374));
    InMux I__10589 (
            .O(N__45408),
            .I(N__45371));
    InMux I__10588 (
            .O(N__45407),
            .I(N__45364));
    InMux I__10587 (
            .O(N__45406),
            .I(N__45364));
    InMux I__10586 (
            .O(N__45405),
            .I(N__45364));
    Span4Mux_v I__10585 (
            .O(N__45402),
            .I(N__45360));
    Span4Mux_v I__10584 (
            .O(N__45399),
            .I(N__45353));
    Span4Mux_v I__10583 (
            .O(N__45396),
            .I(N__45353));
    LocalMux I__10582 (
            .O(N__45383),
            .I(N__45353));
    InMux I__10581 (
            .O(N__45380),
            .I(N__45348));
    InMux I__10580 (
            .O(N__45379),
            .I(N__45348));
    LocalMux I__10579 (
            .O(N__45374),
            .I(N__45345));
    LocalMux I__10578 (
            .O(N__45371),
            .I(N__45340));
    LocalMux I__10577 (
            .O(N__45364),
            .I(N__45340));
    InMux I__10576 (
            .O(N__45363),
            .I(N__45337));
    Span4Mux_h I__10575 (
            .O(N__45360),
            .I(N__45334));
    Span4Mux_h I__10574 (
            .O(N__45353),
            .I(N__45331));
    LocalMux I__10573 (
            .O(N__45348),
            .I(N__45322));
    Span4Mux_v I__10572 (
            .O(N__45345),
            .I(N__45322));
    Span4Mux_h I__10571 (
            .O(N__45340),
            .I(N__45322));
    LocalMux I__10570 (
            .O(N__45337),
            .I(N__45322));
    Odrv4 I__10569 (
            .O(N__45334),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__10568 (
            .O(N__45331),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__10567 (
            .O(N__45322),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__10566 (
            .O(N__45315),
            .I(N__45311));
    InMux I__10565 (
            .O(N__45314),
            .I(N__45308));
    LocalMux I__10564 (
            .O(N__45311),
            .I(N__45305));
    LocalMux I__10563 (
            .O(N__45308),
            .I(N__45302));
    Span4Mux_h I__10562 (
            .O(N__45305),
            .I(N__45299));
    Span4Mux_h I__10561 (
            .O(N__45302),
            .I(N__45296));
    Odrv4 I__10560 (
            .O(N__45299),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__10559 (
            .O(N__45296),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__10558 (
            .O(N__45291),
            .I(N__45288));
    LocalMux I__10557 (
            .O(N__45288),
            .I(N__45285));
    Odrv4 I__10556 (
            .O(N__45285),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    CascadeMux I__10555 (
            .O(N__45282),
            .I(N__45279));
    InMux I__10554 (
            .O(N__45279),
            .I(N__45275));
    InMux I__10553 (
            .O(N__45278),
            .I(N__45272));
    LocalMux I__10552 (
            .O(N__45275),
            .I(N__45269));
    LocalMux I__10551 (
            .O(N__45272),
            .I(N__45266));
    Odrv12 I__10550 (
            .O(N__45269),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__10549 (
            .O(N__45266),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__10548 (
            .O(N__45261),
            .I(N__45258));
    InMux I__10547 (
            .O(N__45258),
            .I(N__45255));
    LocalMux I__10546 (
            .O(N__45255),
            .I(N__45252));
    Odrv12 I__10545 (
            .O(N__45252),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__10544 (
            .O(N__45249),
            .I(N__45245));
    InMux I__10543 (
            .O(N__45248),
            .I(N__45242));
    LocalMux I__10542 (
            .O(N__45245),
            .I(N__45239));
    LocalMux I__10541 (
            .O(N__45242),
            .I(N__45236));
    Odrv12 I__10540 (
            .O(N__45239),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__10539 (
            .O(N__45236),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__10538 (
            .O(N__45231),
            .I(N__45228));
    LocalMux I__10537 (
            .O(N__45228),
            .I(N__45225));
    Odrv4 I__10536 (
            .O(N__45225),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__10535 (
            .O(N__45222),
            .I(N__45218));
    InMux I__10534 (
            .O(N__45221),
            .I(N__45215));
    LocalMux I__10533 (
            .O(N__45218),
            .I(N__45210));
    LocalMux I__10532 (
            .O(N__45215),
            .I(N__45210));
    Odrv4 I__10531 (
            .O(N__45210),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__10530 (
            .O(N__45207),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__10529 (
            .O(N__45204),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__10528 (
            .O(N__45201),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__10527 (
            .O(N__45198),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__10526 (
            .O(N__45195),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__10525 (
            .O(N__45192),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__10524 (
            .O(N__45189),
            .I(N__45185));
    InMux I__10523 (
            .O(N__45188),
            .I(N__45182));
    LocalMux I__10522 (
            .O(N__45185),
            .I(N__45179));
    LocalMux I__10521 (
            .O(N__45182),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__10520 (
            .O(N__45179),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__10519 (
            .O(N__45174),
            .I(N__45171));
    LocalMux I__10518 (
            .O(N__45171),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__10517 (
            .O(N__45168),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__10516 (
            .O(N__45165),
            .I(N__45162));
    LocalMux I__10515 (
            .O(N__45162),
            .I(N__45158));
    InMux I__10514 (
            .O(N__45161),
            .I(N__45155));
    Span4Mux_h I__10513 (
            .O(N__45158),
            .I(N__45152));
    LocalMux I__10512 (
            .O(N__45155),
            .I(N__45149));
    Odrv4 I__10511 (
            .O(N__45152),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__10510 (
            .O(N__45149),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__10509 (
            .O(N__45144),
            .I(N__45141));
    LocalMux I__10508 (
            .O(N__45141),
            .I(N__45138));
    Odrv4 I__10507 (
            .O(N__45138),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    InMux I__10506 (
            .O(N__45135),
            .I(bfn_18_16_0_));
    InMux I__10505 (
            .O(N__45132),
            .I(N__45129));
    LocalMux I__10504 (
            .O(N__45129),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    InMux I__10503 (
            .O(N__45126),
            .I(N__45123));
    LocalMux I__10502 (
            .O(N__45123),
            .I(N__45120));
    Span4Mux_h I__10501 (
            .O(N__45120),
            .I(N__45116));
    InMux I__10500 (
            .O(N__45119),
            .I(N__45113));
    Odrv4 I__10499 (
            .O(N__45116),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__10498 (
            .O(N__45113),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__10497 (
            .O(N__45108),
            .I(N__45105));
    LocalMux I__10496 (
            .O(N__45105),
            .I(N__45102));
    Span4Mux_h I__10495 (
            .O(N__45102),
            .I(N__45099));
    Odrv4 I__10494 (
            .O(N__45099),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    InMux I__10493 (
            .O(N__45096),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__10492 (
            .O(N__45093),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__10491 (
            .O(N__45090),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__10490 (
            .O(N__45087),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__10489 (
            .O(N__45084),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__10488 (
            .O(N__45081),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__10487 (
            .O(N__45078),
            .I(N__45074));
    InMux I__10486 (
            .O(N__45077),
            .I(N__45071));
    LocalMux I__10485 (
            .O(N__45074),
            .I(N__45066));
    LocalMux I__10484 (
            .O(N__45071),
            .I(N__45066));
    Span4Mux_v I__10483 (
            .O(N__45066),
            .I(N__45063));
    Odrv4 I__10482 (
            .O(N__45063),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__10481 (
            .O(N__45060),
            .I(N__45057));
    LocalMux I__10480 (
            .O(N__45057),
            .I(N__45054));
    Span4Mux_h I__10479 (
            .O(N__45054),
            .I(N__45051));
    Odrv4 I__10478 (
            .O(N__45051),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    InMux I__10477 (
            .O(N__45048),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__10476 (
            .O(N__45045),
            .I(N__45041));
    InMux I__10475 (
            .O(N__45044),
            .I(N__45038));
    LocalMux I__10474 (
            .O(N__45041),
            .I(N__45035));
    LocalMux I__10473 (
            .O(N__45038),
            .I(N__45032));
    Span4Mux_v I__10472 (
            .O(N__45035),
            .I(N__45029));
    Span4Mux_v I__10471 (
            .O(N__45032),
            .I(N__45026));
    Odrv4 I__10470 (
            .O(N__45029),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__10469 (
            .O(N__45026),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__10468 (
            .O(N__45021),
            .I(N__45018));
    LocalMux I__10467 (
            .O(N__45018),
            .I(N__45015));
    Span4Mux_h I__10466 (
            .O(N__45015),
            .I(N__45012));
    Odrv4 I__10465 (
            .O(N__45012),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    InMux I__10464 (
            .O(N__45009),
            .I(bfn_18_15_0_));
    InMux I__10463 (
            .O(N__45006),
            .I(N__45002));
    InMux I__10462 (
            .O(N__45005),
            .I(N__44999));
    LocalMux I__10461 (
            .O(N__45002),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__10460 (
            .O(N__44999),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__10459 (
            .O(N__44994),
            .I(N__44991));
    InMux I__10458 (
            .O(N__44991),
            .I(N__44988));
    LocalMux I__10457 (
            .O(N__44988),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ));
    InMux I__10456 (
            .O(N__44985),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__10455 (
            .O(N__44982),
            .I(N__44978));
    InMux I__10454 (
            .O(N__44981),
            .I(N__44975));
    LocalMux I__10453 (
            .O(N__44978),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__10452 (
            .O(N__44975),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__10451 (
            .O(N__44970),
            .I(N__44967));
    LocalMux I__10450 (
            .O(N__44967),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ));
    InMux I__10449 (
            .O(N__44964),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__10448 (
            .O(N__44961),
            .I(N__44957));
    InMux I__10447 (
            .O(N__44960),
            .I(N__44954));
    LocalMux I__10446 (
            .O(N__44957),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__10445 (
            .O(N__44954),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__10444 (
            .O(N__44949),
            .I(N__44946));
    InMux I__10443 (
            .O(N__44946),
            .I(N__44943));
    LocalMux I__10442 (
            .O(N__44943),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__10441 (
            .O(N__44940),
            .I(bfn_18_13_0_));
    InMux I__10440 (
            .O(N__44937),
            .I(N__44933));
    InMux I__10439 (
            .O(N__44936),
            .I(N__44930));
    LocalMux I__10438 (
            .O(N__44933),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__10437 (
            .O(N__44930),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__10436 (
            .O(N__44925),
            .I(N__44922));
    LocalMux I__10435 (
            .O(N__44922),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__10434 (
            .O(N__44919),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__10433 (
            .O(N__44916),
            .I(N__44912));
    InMux I__10432 (
            .O(N__44915),
            .I(N__44909));
    LocalMux I__10431 (
            .O(N__44912),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__10430 (
            .O(N__44909),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__10429 (
            .O(N__44904),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ));
    CascadeMux I__10428 (
            .O(N__44901),
            .I(N__44898));
    InMux I__10427 (
            .O(N__44898),
            .I(N__44895));
    LocalMux I__10426 (
            .O(N__44895),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ));
    InMux I__10425 (
            .O(N__44892),
            .I(N__44868));
    InMux I__10424 (
            .O(N__44891),
            .I(N__44868));
    InMux I__10423 (
            .O(N__44890),
            .I(N__44851));
    InMux I__10422 (
            .O(N__44889),
            .I(N__44851));
    InMux I__10421 (
            .O(N__44888),
            .I(N__44851));
    InMux I__10420 (
            .O(N__44887),
            .I(N__44851));
    InMux I__10419 (
            .O(N__44886),
            .I(N__44851));
    InMux I__10418 (
            .O(N__44885),
            .I(N__44851));
    InMux I__10417 (
            .O(N__44884),
            .I(N__44851));
    InMux I__10416 (
            .O(N__44883),
            .I(N__44851));
    InMux I__10415 (
            .O(N__44882),
            .I(N__44834));
    InMux I__10414 (
            .O(N__44881),
            .I(N__44834));
    InMux I__10413 (
            .O(N__44880),
            .I(N__44834));
    InMux I__10412 (
            .O(N__44879),
            .I(N__44834));
    InMux I__10411 (
            .O(N__44878),
            .I(N__44834));
    InMux I__10410 (
            .O(N__44877),
            .I(N__44834));
    InMux I__10409 (
            .O(N__44876),
            .I(N__44834));
    InMux I__10408 (
            .O(N__44875),
            .I(N__44834));
    InMux I__10407 (
            .O(N__44874),
            .I(N__44831));
    InMux I__10406 (
            .O(N__44873),
            .I(N__44828));
    LocalMux I__10405 (
            .O(N__44868),
            .I(N__44823));
    LocalMux I__10404 (
            .O(N__44851),
            .I(N__44823));
    LocalMux I__10403 (
            .O(N__44834),
            .I(N__44814));
    LocalMux I__10402 (
            .O(N__44831),
            .I(N__44814));
    LocalMux I__10401 (
            .O(N__44828),
            .I(N__44811));
    Span4Mux_h I__10400 (
            .O(N__44823),
            .I(N__44808));
    InMux I__10399 (
            .O(N__44822),
            .I(N__44805));
    InMux I__10398 (
            .O(N__44821),
            .I(N__44802));
    InMux I__10397 (
            .O(N__44820),
            .I(N__44797));
    InMux I__10396 (
            .O(N__44819),
            .I(N__44797));
    Span4Mux_h I__10395 (
            .O(N__44814),
            .I(N__44794));
    Span4Mux_v I__10394 (
            .O(N__44811),
            .I(N__44787));
    Span4Mux_h I__10393 (
            .O(N__44808),
            .I(N__44787));
    LocalMux I__10392 (
            .O(N__44805),
            .I(N__44787));
    LocalMux I__10391 (
            .O(N__44802),
            .I(N__44784));
    LocalMux I__10390 (
            .O(N__44797),
            .I(N__44779));
    Span4Mux_v I__10389 (
            .O(N__44794),
            .I(N__44779));
    Odrv4 I__10388 (
            .O(N__44787),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv12 I__10387 (
            .O(N__44784),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__10386 (
            .O(N__44779),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__10385 (
            .O(N__44772),
            .I(N__44760));
    InMux I__10384 (
            .O(N__44771),
            .I(N__44733));
    InMux I__10383 (
            .O(N__44770),
            .I(N__44733));
    InMux I__10382 (
            .O(N__44769),
            .I(N__44733));
    InMux I__10381 (
            .O(N__44768),
            .I(N__44733));
    InMux I__10380 (
            .O(N__44767),
            .I(N__44733));
    InMux I__10379 (
            .O(N__44766),
            .I(N__44733));
    InMux I__10378 (
            .O(N__44765),
            .I(N__44733));
    InMux I__10377 (
            .O(N__44764),
            .I(N__44733));
    InMux I__10376 (
            .O(N__44763),
            .I(N__44730));
    InMux I__10375 (
            .O(N__44760),
            .I(N__44726));
    InMux I__10374 (
            .O(N__44759),
            .I(N__44709));
    InMux I__10373 (
            .O(N__44758),
            .I(N__44709));
    InMux I__10372 (
            .O(N__44757),
            .I(N__44709));
    InMux I__10371 (
            .O(N__44756),
            .I(N__44709));
    InMux I__10370 (
            .O(N__44755),
            .I(N__44709));
    InMux I__10369 (
            .O(N__44754),
            .I(N__44709));
    InMux I__10368 (
            .O(N__44753),
            .I(N__44709));
    InMux I__10367 (
            .O(N__44752),
            .I(N__44709));
    InMux I__10366 (
            .O(N__44751),
            .I(N__44702));
    InMux I__10365 (
            .O(N__44750),
            .I(N__44702));
    LocalMux I__10364 (
            .O(N__44733),
            .I(N__44697));
    LocalMux I__10363 (
            .O(N__44730),
            .I(N__44697));
    CascadeMux I__10362 (
            .O(N__44729),
            .I(N__44693));
    LocalMux I__10361 (
            .O(N__44726),
            .I(N__44690));
    LocalMux I__10360 (
            .O(N__44709),
            .I(N__44687));
    InMux I__10359 (
            .O(N__44708),
            .I(N__44684));
    InMux I__10358 (
            .O(N__44707),
            .I(N__44681));
    LocalMux I__10357 (
            .O(N__44702),
            .I(N__44676));
    Span4Mux_h I__10356 (
            .O(N__44697),
            .I(N__44676));
    InMux I__10355 (
            .O(N__44696),
            .I(N__44671));
    InMux I__10354 (
            .O(N__44693),
            .I(N__44671));
    Span4Mux_v I__10353 (
            .O(N__44690),
            .I(N__44664));
    Span4Mux_h I__10352 (
            .O(N__44687),
            .I(N__44664));
    LocalMux I__10351 (
            .O(N__44684),
            .I(N__44664));
    LocalMux I__10350 (
            .O(N__44681),
            .I(N__44661));
    Span4Mux_v I__10349 (
            .O(N__44676),
            .I(N__44658));
    LocalMux I__10348 (
            .O(N__44671),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__10347 (
            .O(N__44664),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv12 I__10346 (
            .O(N__44661),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__10345 (
            .O(N__44658),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    InMux I__10344 (
            .O(N__44649),
            .I(N__44644));
    InMux I__10343 (
            .O(N__44648),
            .I(N__44638));
    InMux I__10342 (
            .O(N__44647),
            .I(N__44638));
    LocalMux I__10341 (
            .O(N__44644),
            .I(N__44635));
    InMux I__10340 (
            .O(N__44643),
            .I(N__44632));
    LocalMux I__10339 (
            .O(N__44638),
            .I(N__44629));
    Odrv12 I__10338 (
            .O(N__44635),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    LocalMux I__10337 (
            .O(N__44632),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    Odrv4 I__10336 (
            .O(N__44629),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    InMux I__10335 (
            .O(N__44622),
            .I(N__44615));
    InMux I__10334 (
            .O(N__44621),
            .I(N__44615));
    InMux I__10333 (
            .O(N__44620),
            .I(N__44612));
    LocalMux I__10332 (
            .O(N__44615),
            .I(N__44608));
    LocalMux I__10331 (
            .O(N__44612),
            .I(N__44604));
    InMux I__10330 (
            .O(N__44611),
            .I(N__44601));
    Span4Mux_h I__10329 (
            .O(N__44608),
            .I(N__44598));
    InMux I__10328 (
            .O(N__44607),
            .I(N__44595));
    Span4Mux_h I__10327 (
            .O(N__44604),
            .I(N__44590));
    LocalMux I__10326 (
            .O(N__44601),
            .I(N__44590));
    Odrv4 I__10325 (
            .O(N__44598),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__10324 (
            .O(N__44595),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__10323 (
            .O(N__44590),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__10322 (
            .O(N__44583),
            .I(N__44580));
    LocalMux I__10321 (
            .O(N__44580),
            .I(N__44577));
    Odrv4 I__10320 (
            .O(N__44577),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ));
    InMux I__10319 (
            .O(N__44574),
            .I(N__44570));
    InMux I__10318 (
            .O(N__44573),
            .I(N__44567));
    LocalMux I__10317 (
            .O(N__44570),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__10316 (
            .O(N__44567),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__10315 (
            .O(N__44562),
            .I(N__44559));
    InMux I__10314 (
            .O(N__44559),
            .I(N__44556));
    LocalMux I__10313 (
            .O(N__44556),
            .I(N__44553));
    Odrv4 I__10312 (
            .O(N__44553),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ));
    InMux I__10311 (
            .O(N__44550),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__10310 (
            .O(N__44547),
            .I(N__44543));
    InMux I__10309 (
            .O(N__44546),
            .I(N__44540));
    LocalMux I__10308 (
            .O(N__44543),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__10307 (
            .O(N__44540),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__10306 (
            .O(N__44535),
            .I(N__44532));
    LocalMux I__10305 (
            .O(N__44532),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ));
    InMux I__10304 (
            .O(N__44529),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__10303 (
            .O(N__44526),
            .I(N__44522));
    InMux I__10302 (
            .O(N__44525),
            .I(N__44519));
    LocalMux I__10301 (
            .O(N__44522),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__10300 (
            .O(N__44519),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__10299 (
            .O(N__44514),
            .I(N__44511));
    LocalMux I__10298 (
            .O(N__44511),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ));
    InMux I__10297 (
            .O(N__44508),
            .I(bfn_18_12_0_));
    InMux I__10296 (
            .O(N__44505),
            .I(N__44501));
    InMux I__10295 (
            .O(N__44504),
            .I(N__44498));
    LocalMux I__10294 (
            .O(N__44501),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__10293 (
            .O(N__44498),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__10292 (
            .O(N__44493),
            .I(N__44490));
    LocalMux I__10291 (
            .O(N__44490),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__10290 (
            .O(N__44487),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__10289 (
            .O(N__44484),
            .I(N__44481));
    LocalMux I__10288 (
            .O(N__44481),
            .I(N__44477));
    InMux I__10287 (
            .O(N__44480),
            .I(N__44474));
    Odrv12 I__10286 (
            .O(N__44477),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__10285 (
            .O(N__44474),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__10284 (
            .O(N__44469),
            .I(N__44466));
    InMux I__10283 (
            .O(N__44466),
            .I(N__44463));
    LocalMux I__10282 (
            .O(N__44463),
            .I(N__44460));
    Odrv4 I__10281 (
            .O(N__44460),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ));
    InMux I__10280 (
            .O(N__44457),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__10279 (
            .O(N__44454),
            .I(N__44450));
    InMux I__10278 (
            .O(N__44453),
            .I(N__44447));
    LocalMux I__10277 (
            .O(N__44450),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__10276 (
            .O(N__44447),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__10275 (
            .O(N__44442),
            .I(N__44439));
    InMux I__10274 (
            .O(N__44439),
            .I(N__44436));
    LocalMux I__10273 (
            .O(N__44436),
            .I(N__44433));
    Odrv4 I__10272 (
            .O(N__44433),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__10271 (
            .O(N__44430),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__10270 (
            .O(N__44427),
            .I(N__44424));
    LocalMux I__10269 (
            .O(N__44424),
            .I(N__44420));
    InMux I__10268 (
            .O(N__44423),
            .I(N__44417));
    Span4Mux_h I__10267 (
            .O(N__44420),
            .I(N__44412));
    LocalMux I__10266 (
            .O(N__44417),
            .I(N__44412));
    Span4Mux_h I__10265 (
            .O(N__44412),
            .I(N__44409));
    Odrv4 I__10264 (
            .O(N__44409),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__10263 (
            .O(N__44406),
            .I(N__44403));
    LocalMux I__10262 (
            .O(N__44403),
            .I(N__44400));
    Span4Mux_v I__10261 (
            .O(N__44400),
            .I(N__44397));
    Odrv4 I__10260 (
            .O(N__44397),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ));
    InMux I__10259 (
            .O(N__44394),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__10258 (
            .O(N__44391),
            .I(N__44387));
    InMux I__10257 (
            .O(N__44390),
            .I(N__44384));
    LocalMux I__10256 (
            .O(N__44387),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__10255 (
            .O(N__44384),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__10254 (
            .O(N__44379),
            .I(N__44376));
    InMux I__10253 (
            .O(N__44376),
            .I(N__44373));
    LocalMux I__10252 (
            .O(N__44373),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ));
    InMux I__10251 (
            .O(N__44370),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ));
    CascadeMux I__10250 (
            .O(N__44367),
            .I(N__44363));
    InMux I__10249 (
            .O(N__44366),
            .I(N__44360));
    InMux I__10248 (
            .O(N__44363),
            .I(N__44357));
    LocalMux I__10247 (
            .O(N__44360),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__10246 (
            .O(N__44357),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__10245 (
            .O(N__44352),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__10244 (
            .O(N__44349),
            .I(N__44311));
    InMux I__10243 (
            .O(N__44348),
            .I(N__44311));
    InMux I__10242 (
            .O(N__44347),
            .I(N__44311));
    InMux I__10241 (
            .O(N__44346),
            .I(N__44311));
    InMux I__10240 (
            .O(N__44345),
            .I(N__44302));
    InMux I__10239 (
            .O(N__44344),
            .I(N__44302));
    InMux I__10238 (
            .O(N__44343),
            .I(N__44302));
    InMux I__10237 (
            .O(N__44342),
            .I(N__44302));
    InMux I__10236 (
            .O(N__44341),
            .I(N__44293));
    InMux I__10235 (
            .O(N__44340),
            .I(N__44293));
    InMux I__10234 (
            .O(N__44339),
            .I(N__44293));
    InMux I__10233 (
            .O(N__44338),
            .I(N__44293));
    InMux I__10232 (
            .O(N__44337),
            .I(N__44284));
    InMux I__10231 (
            .O(N__44336),
            .I(N__44284));
    InMux I__10230 (
            .O(N__44335),
            .I(N__44284));
    InMux I__10229 (
            .O(N__44334),
            .I(N__44284));
    InMux I__10228 (
            .O(N__44333),
            .I(N__44275));
    InMux I__10227 (
            .O(N__44332),
            .I(N__44275));
    InMux I__10226 (
            .O(N__44331),
            .I(N__44275));
    InMux I__10225 (
            .O(N__44330),
            .I(N__44275));
    InMux I__10224 (
            .O(N__44329),
            .I(N__44270));
    InMux I__10223 (
            .O(N__44328),
            .I(N__44270));
    InMux I__10222 (
            .O(N__44327),
            .I(N__44261));
    InMux I__10221 (
            .O(N__44326),
            .I(N__44261));
    InMux I__10220 (
            .O(N__44325),
            .I(N__44261));
    InMux I__10219 (
            .O(N__44324),
            .I(N__44261));
    InMux I__10218 (
            .O(N__44323),
            .I(N__44252));
    InMux I__10217 (
            .O(N__44322),
            .I(N__44252));
    InMux I__10216 (
            .O(N__44321),
            .I(N__44252));
    InMux I__10215 (
            .O(N__44320),
            .I(N__44252));
    LocalMux I__10214 (
            .O(N__44311),
            .I(N__44243));
    LocalMux I__10213 (
            .O(N__44302),
            .I(N__44243));
    LocalMux I__10212 (
            .O(N__44293),
            .I(N__44243));
    LocalMux I__10211 (
            .O(N__44284),
            .I(N__44243));
    LocalMux I__10210 (
            .O(N__44275),
            .I(N__44236));
    LocalMux I__10209 (
            .O(N__44270),
            .I(N__44236));
    LocalMux I__10208 (
            .O(N__44261),
            .I(N__44236));
    LocalMux I__10207 (
            .O(N__44252),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__10206 (
            .O(N__44243),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv12 I__10205 (
            .O(N__44236),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__10204 (
            .O(N__44229),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CascadeMux I__10203 (
            .O(N__44226),
            .I(N__44222));
    InMux I__10202 (
            .O(N__44225),
            .I(N__44219));
    InMux I__10201 (
            .O(N__44222),
            .I(N__44216));
    LocalMux I__10200 (
            .O(N__44219),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__10199 (
            .O(N__44216),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CEMux I__10198 (
            .O(N__44211),
            .I(N__44208));
    LocalMux I__10197 (
            .O(N__44208),
            .I(N__44202));
    CEMux I__10196 (
            .O(N__44207),
            .I(N__44199));
    CEMux I__10195 (
            .O(N__44206),
            .I(N__44196));
    CEMux I__10194 (
            .O(N__44205),
            .I(N__44193));
    Span4Mux_v I__10193 (
            .O(N__44202),
            .I(N__44188));
    LocalMux I__10192 (
            .O(N__44199),
            .I(N__44188));
    LocalMux I__10191 (
            .O(N__44196),
            .I(N__44183));
    LocalMux I__10190 (
            .O(N__44193),
            .I(N__44183));
    Span4Mux_v I__10189 (
            .O(N__44188),
            .I(N__44178));
    Span4Mux_v I__10188 (
            .O(N__44183),
            .I(N__44178));
    Odrv4 I__10187 (
            .O(N__44178),
            .I(\delay_measurement_inst.delay_hc_timer.N_336_i ));
    InMux I__10186 (
            .O(N__44175),
            .I(N__44172));
    LocalMux I__10185 (
            .O(N__44172),
            .I(N__44169));
    Span4Mux_h I__10184 (
            .O(N__44169),
            .I(N__44166));
    Odrv4 I__10183 (
            .O(N__44166),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    CascadeMux I__10182 (
            .O(N__44163),
            .I(N__44160));
    InMux I__10181 (
            .O(N__44160),
            .I(N__44157));
    LocalMux I__10180 (
            .O(N__44157),
            .I(N__44153));
    InMux I__10179 (
            .O(N__44156),
            .I(N__44149));
    Span4Mux_h I__10178 (
            .O(N__44153),
            .I(N__44146));
    InMux I__10177 (
            .O(N__44152),
            .I(N__44143));
    LocalMux I__10176 (
            .O(N__44149),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__10175 (
            .O(N__44146),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__10174 (
            .O(N__44143),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__10173 (
            .O(N__44136),
            .I(N__44132));
    InMux I__10172 (
            .O(N__44135),
            .I(N__44129));
    LocalMux I__10171 (
            .O(N__44132),
            .I(N__44126));
    LocalMux I__10170 (
            .O(N__44129),
            .I(N__44123));
    Odrv4 I__10169 (
            .O(N__44126),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__10168 (
            .O(N__44123),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__10167 (
            .O(N__44118),
            .I(N__44115));
    LocalMux I__10166 (
            .O(N__44115),
            .I(N__44112));
    Span4Mux_h I__10165 (
            .O(N__44112),
            .I(N__44109));
    Odrv4 I__10164 (
            .O(N__44109),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ));
    InMux I__10163 (
            .O(N__44106),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ));
    CascadeMux I__10162 (
            .O(N__44103),
            .I(N__44100));
    InMux I__10161 (
            .O(N__44100),
            .I(N__44096));
    InMux I__10160 (
            .O(N__44099),
            .I(N__44093));
    LocalMux I__10159 (
            .O(N__44096),
            .I(N__44090));
    LocalMux I__10158 (
            .O(N__44093),
            .I(N__44087));
    Odrv4 I__10157 (
            .O(N__44090),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__10156 (
            .O(N__44087),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__10155 (
            .O(N__44082),
            .I(N__44079));
    InMux I__10154 (
            .O(N__44079),
            .I(N__44076));
    LocalMux I__10153 (
            .O(N__44076),
            .I(N__44073));
    Span4Mux_v I__10152 (
            .O(N__44073),
            .I(N__44070));
    Odrv4 I__10151 (
            .O(N__44070),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ));
    InMux I__10150 (
            .O(N__44067),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__10149 (
            .O(N__44064),
            .I(N__44060));
    InMux I__10148 (
            .O(N__44063),
            .I(N__44057));
    LocalMux I__10147 (
            .O(N__44060),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__10146 (
            .O(N__44057),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__10145 (
            .O(N__44052),
            .I(N__44049));
    LocalMux I__10144 (
            .O(N__44049),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ));
    InMux I__10143 (
            .O(N__44046),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__10142 (
            .O(N__44043),
            .I(N__44039));
    InMux I__10141 (
            .O(N__44042),
            .I(N__44036));
    LocalMux I__10140 (
            .O(N__44039),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__10139 (
            .O(N__44036),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__10138 (
            .O(N__44031),
            .I(N__44028));
    InMux I__10137 (
            .O(N__44028),
            .I(N__44025));
    LocalMux I__10136 (
            .O(N__44025),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ));
    InMux I__10135 (
            .O(N__44022),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__10134 (
            .O(N__44019),
            .I(N__44015));
    InMux I__10133 (
            .O(N__44018),
            .I(N__44012));
    LocalMux I__10132 (
            .O(N__44015),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__10131 (
            .O(N__44012),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__10130 (
            .O(N__44007),
            .I(N__44004));
    LocalMux I__10129 (
            .O(N__44004),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ));
    InMux I__10128 (
            .O(N__44001),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ));
    CascadeMux I__10127 (
            .O(N__43998),
            .I(N__43993));
    InMux I__10126 (
            .O(N__43997),
            .I(N__43990));
    InMux I__10125 (
            .O(N__43996),
            .I(N__43987));
    InMux I__10124 (
            .O(N__43993),
            .I(N__43984));
    LocalMux I__10123 (
            .O(N__43990),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__10122 (
            .O(N__43987),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__10121 (
            .O(N__43984),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__10120 (
            .O(N__43977),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__10119 (
            .O(N__43974),
            .I(N__43969));
    InMux I__10118 (
            .O(N__43973),
            .I(N__43966));
    InMux I__10117 (
            .O(N__43972),
            .I(N__43963));
    InMux I__10116 (
            .O(N__43969),
            .I(N__43960));
    LocalMux I__10115 (
            .O(N__43966),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__10114 (
            .O(N__43963),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__10113 (
            .O(N__43960),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__10112 (
            .O(N__43953),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    CascadeMux I__10111 (
            .O(N__43950),
            .I(N__43945));
    InMux I__10110 (
            .O(N__43949),
            .I(N__43942));
    InMux I__10109 (
            .O(N__43948),
            .I(N__43939));
    InMux I__10108 (
            .O(N__43945),
            .I(N__43936));
    LocalMux I__10107 (
            .O(N__43942),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__10106 (
            .O(N__43939),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__10105 (
            .O(N__43936),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__10104 (
            .O(N__43929),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    CascadeMux I__10103 (
            .O(N__43926),
            .I(N__43921));
    InMux I__10102 (
            .O(N__43925),
            .I(N__43918));
    InMux I__10101 (
            .O(N__43924),
            .I(N__43915));
    InMux I__10100 (
            .O(N__43921),
            .I(N__43912));
    LocalMux I__10099 (
            .O(N__43918),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__10098 (
            .O(N__43915),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__10097 (
            .O(N__43912),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__10096 (
            .O(N__43905),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__10095 (
            .O(N__43902),
            .I(N__43897));
    InMux I__10094 (
            .O(N__43901),
            .I(N__43894));
    InMux I__10093 (
            .O(N__43900),
            .I(N__43891));
    InMux I__10092 (
            .O(N__43897),
            .I(N__43888));
    LocalMux I__10091 (
            .O(N__43894),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__10090 (
            .O(N__43891),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__10089 (
            .O(N__43888),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__10088 (
            .O(N__43881),
            .I(bfn_18_10_0_));
    CascadeMux I__10087 (
            .O(N__43878),
            .I(N__43873));
    InMux I__10086 (
            .O(N__43877),
            .I(N__43870));
    InMux I__10085 (
            .O(N__43876),
            .I(N__43867));
    InMux I__10084 (
            .O(N__43873),
            .I(N__43864));
    LocalMux I__10083 (
            .O(N__43870),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__10082 (
            .O(N__43867),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__10081 (
            .O(N__43864),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__10080 (
            .O(N__43857),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__10079 (
            .O(N__43854),
            .I(N__43849));
    InMux I__10078 (
            .O(N__43853),
            .I(N__43846));
    InMux I__10077 (
            .O(N__43852),
            .I(N__43843));
    InMux I__10076 (
            .O(N__43849),
            .I(N__43840));
    LocalMux I__10075 (
            .O(N__43846),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__10074 (
            .O(N__43843),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__10073 (
            .O(N__43840),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__10072 (
            .O(N__43833),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__10071 (
            .O(N__43830),
            .I(N__43825));
    InMux I__10070 (
            .O(N__43829),
            .I(N__43822));
    InMux I__10069 (
            .O(N__43828),
            .I(N__43819));
    InMux I__10068 (
            .O(N__43825),
            .I(N__43816));
    LocalMux I__10067 (
            .O(N__43822),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__10066 (
            .O(N__43819),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__10065 (
            .O(N__43816),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__10064 (
            .O(N__43809),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    CascadeMux I__10063 (
            .O(N__43806),
            .I(N__43801));
    InMux I__10062 (
            .O(N__43805),
            .I(N__43798));
    InMux I__10061 (
            .O(N__43804),
            .I(N__43795));
    InMux I__10060 (
            .O(N__43801),
            .I(N__43792));
    LocalMux I__10059 (
            .O(N__43798),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__10058 (
            .O(N__43795),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__10057 (
            .O(N__43792),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__10056 (
            .O(N__43785),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    CascadeMux I__10055 (
            .O(N__43782),
            .I(N__43777));
    InMux I__10054 (
            .O(N__43781),
            .I(N__43774));
    InMux I__10053 (
            .O(N__43780),
            .I(N__43771));
    InMux I__10052 (
            .O(N__43777),
            .I(N__43768));
    LocalMux I__10051 (
            .O(N__43774),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__10050 (
            .O(N__43771),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__10049 (
            .O(N__43768),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__10048 (
            .O(N__43761),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    CascadeMux I__10047 (
            .O(N__43758),
            .I(N__43753));
    InMux I__10046 (
            .O(N__43757),
            .I(N__43750));
    InMux I__10045 (
            .O(N__43756),
            .I(N__43747));
    InMux I__10044 (
            .O(N__43753),
            .I(N__43744));
    LocalMux I__10043 (
            .O(N__43750),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__10042 (
            .O(N__43747),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__10041 (
            .O(N__43744),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__10040 (
            .O(N__43737),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    CascadeMux I__10039 (
            .O(N__43734),
            .I(N__43729));
    InMux I__10038 (
            .O(N__43733),
            .I(N__43726));
    InMux I__10037 (
            .O(N__43732),
            .I(N__43723));
    InMux I__10036 (
            .O(N__43729),
            .I(N__43720));
    LocalMux I__10035 (
            .O(N__43726),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__10034 (
            .O(N__43723),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__10033 (
            .O(N__43720),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__10032 (
            .O(N__43713),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__10031 (
            .O(N__43710),
            .I(N__43705));
    InMux I__10030 (
            .O(N__43709),
            .I(N__43702));
    InMux I__10029 (
            .O(N__43708),
            .I(N__43699));
    InMux I__10028 (
            .O(N__43705),
            .I(N__43696));
    LocalMux I__10027 (
            .O(N__43702),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__10026 (
            .O(N__43699),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__10025 (
            .O(N__43696),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__10024 (
            .O(N__43689),
            .I(bfn_18_9_0_));
    CascadeMux I__10023 (
            .O(N__43686),
            .I(N__43681));
    InMux I__10022 (
            .O(N__43685),
            .I(N__43678));
    InMux I__10021 (
            .O(N__43684),
            .I(N__43675));
    InMux I__10020 (
            .O(N__43681),
            .I(N__43672));
    LocalMux I__10019 (
            .O(N__43678),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__10018 (
            .O(N__43675),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__10017 (
            .O(N__43672),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__10016 (
            .O(N__43665),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__10015 (
            .O(N__43662),
            .I(N__43657));
    InMux I__10014 (
            .O(N__43661),
            .I(N__43654));
    InMux I__10013 (
            .O(N__43660),
            .I(N__43651));
    InMux I__10012 (
            .O(N__43657),
            .I(N__43648));
    LocalMux I__10011 (
            .O(N__43654),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__10010 (
            .O(N__43651),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__10009 (
            .O(N__43648),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__10008 (
            .O(N__43641),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__10007 (
            .O(N__43638),
            .I(N__43633));
    InMux I__10006 (
            .O(N__43637),
            .I(N__43630));
    InMux I__10005 (
            .O(N__43636),
            .I(N__43627));
    InMux I__10004 (
            .O(N__43633),
            .I(N__43624));
    LocalMux I__10003 (
            .O(N__43630),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__10002 (
            .O(N__43627),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__10001 (
            .O(N__43624),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__10000 (
            .O(N__43617),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    CascadeMux I__9999 (
            .O(N__43614),
            .I(N__43609));
    InMux I__9998 (
            .O(N__43613),
            .I(N__43606));
    InMux I__9997 (
            .O(N__43612),
            .I(N__43603));
    InMux I__9996 (
            .O(N__43609),
            .I(N__43600));
    LocalMux I__9995 (
            .O(N__43606),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__9994 (
            .O(N__43603),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__9993 (
            .O(N__43600),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__9992 (
            .O(N__43593),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__9991 (
            .O(N__43590),
            .I(N__43585));
    InMux I__9990 (
            .O(N__43589),
            .I(N__43582));
    InMux I__9989 (
            .O(N__43588),
            .I(N__43579));
    InMux I__9988 (
            .O(N__43585),
            .I(N__43576));
    LocalMux I__9987 (
            .O(N__43582),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__9986 (
            .O(N__43579),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__9985 (
            .O(N__43576),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__9984 (
            .O(N__43569),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__9983 (
            .O(N__43566),
            .I(N__43561));
    InMux I__9982 (
            .O(N__43565),
            .I(N__43558));
    InMux I__9981 (
            .O(N__43564),
            .I(N__43555));
    InMux I__9980 (
            .O(N__43561),
            .I(N__43552));
    LocalMux I__9979 (
            .O(N__43558),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__9978 (
            .O(N__43555),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__9977 (
            .O(N__43552),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__9976 (
            .O(N__43545),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    CascadeMux I__9975 (
            .O(N__43542),
            .I(N__43537));
    InMux I__9974 (
            .O(N__43541),
            .I(N__43534));
    InMux I__9973 (
            .O(N__43540),
            .I(N__43531));
    InMux I__9972 (
            .O(N__43537),
            .I(N__43528));
    LocalMux I__9971 (
            .O(N__43534),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__9970 (
            .O(N__43531),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__9969 (
            .O(N__43528),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__9968 (
            .O(N__43521),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    CascadeMux I__9967 (
            .O(N__43518),
            .I(N__43513));
    InMux I__9966 (
            .O(N__43517),
            .I(N__43510));
    InMux I__9965 (
            .O(N__43516),
            .I(N__43507));
    InMux I__9964 (
            .O(N__43513),
            .I(N__43504));
    LocalMux I__9963 (
            .O(N__43510),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__9962 (
            .O(N__43507),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__9961 (
            .O(N__43504),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__9960 (
            .O(N__43497),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__9959 (
            .O(N__43494),
            .I(N__43489));
    InMux I__9958 (
            .O(N__43493),
            .I(N__43486));
    InMux I__9957 (
            .O(N__43492),
            .I(N__43483));
    InMux I__9956 (
            .O(N__43489),
            .I(N__43480));
    LocalMux I__9955 (
            .O(N__43486),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__9954 (
            .O(N__43483),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__9953 (
            .O(N__43480),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__9952 (
            .O(N__43473),
            .I(bfn_18_8_0_));
    CascadeMux I__9951 (
            .O(N__43470),
            .I(N__43465));
    InMux I__9950 (
            .O(N__43469),
            .I(N__43462));
    InMux I__9949 (
            .O(N__43468),
            .I(N__43459));
    InMux I__9948 (
            .O(N__43465),
            .I(N__43456));
    LocalMux I__9947 (
            .O(N__43462),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__9946 (
            .O(N__43459),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__9945 (
            .O(N__43456),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__9944 (
            .O(N__43449),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    CascadeMux I__9943 (
            .O(N__43446),
            .I(N__43441));
    InMux I__9942 (
            .O(N__43445),
            .I(N__43438));
    InMux I__9941 (
            .O(N__43444),
            .I(N__43435));
    InMux I__9940 (
            .O(N__43441),
            .I(N__43432));
    LocalMux I__9939 (
            .O(N__43438),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__9938 (
            .O(N__43435),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__9937 (
            .O(N__43432),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__9936 (
            .O(N__43425),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    CascadeMux I__9935 (
            .O(N__43422),
            .I(N__43417));
    InMux I__9934 (
            .O(N__43421),
            .I(N__43414));
    InMux I__9933 (
            .O(N__43420),
            .I(N__43411));
    InMux I__9932 (
            .O(N__43417),
            .I(N__43408));
    LocalMux I__9931 (
            .O(N__43414),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__9930 (
            .O(N__43411),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__9929 (
            .O(N__43408),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__9928 (
            .O(N__43401),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    CascadeMux I__9927 (
            .O(N__43398),
            .I(N__43395));
    InMux I__9926 (
            .O(N__43395),
            .I(N__43392));
    LocalMux I__9925 (
            .O(N__43392),
            .I(N__43389));
    Odrv4 I__9924 (
            .O(N__43389),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ));
    CEMux I__9923 (
            .O(N__43386),
            .I(N__43381));
    CEMux I__9922 (
            .O(N__43385),
            .I(N__43377));
    CEMux I__9921 (
            .O(N__43384),
            .I(N__43374));
    LocalMux I__9920 (
            .O(N__43381),
            .I(N__43371));
    CEMux I__9919 (
            .O(N__43380),
            .I(N__43368));
    LocalMux I__9918 (
            .O(N__43377),
            .I(N__43365));
    LocalMux I__9917 (
            .O(N__43374),
            .I(N__43362));
    Span4Mux_v I__9916 (
            .O(N__43371),
            .I(N__43357));
    LocalMux I__9915 (
            .O(N__43368),
            .I(N__43357));
    Span4Mux_v I__9914 (
            .O(N__43365),
            .I(N__43352));
    Span4Mux_v I__9913 (
            .O(N__43362),
            .I(N__43352));
    Span4Mux_v I__9912 (
            .O(N__43357),
            .I(N__43349));
    Odrv4 I__9911 (
            .O(N__43352),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__9910 (
            .O(N__43349),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    CascadeMux I__9909 (
            .O(N__43344),
            .I(N__43336));
    CascadeMux I__9908 (
            .O(N__43343),
            .I(N__43333));
    InMux I__9907 (
            .O(N__43342),
            .I(N__43319));
    InMux I__9906 (
            .O(N__43341),
            .I(N__43319));
    InMux I__9905 (
            .O(N__43340),
            .I(N__43319));
    InMux I__9904 (
            .O(N__43339),
            .I(N__43319));
    InMux I__9903 (
            .O(N__43336),
            .I(N__43306));
    InMux I__9902 (
            .O(N__43333),
            .I(N__43306));
    InMux I__9901 (
            .O(N__43332),
            .I(N__43306));
    InMux I__9900 (
            .O(N__43331),
            .I(N__43306));
    InMux I__9899 (
            .O(N__43330),
            .I(N__43306));
    InMux I__9898 (
            .O(N__43329),
            .I(N__43306));
    InMux I__9897 (
            .O(N__43328),
            .I(N__43303));
    LocalMux I__9896 (
            .O(N__43319),
            .I(N__43296));
    LocalMux I__9895 (
            .O(N__43306),
            .I(N__43293));
    LocalMux I__9894 (
            .O(N__43303),
            .I(N__43290));
    InMux I__9893 (
            .O(N__43302),
            .I(N__43287));
    InMux I__9892 (
            .O(N__43301),
            .I(N__43282));
    InMux I__9891 (
            .O(N__43300),
            .I(N__43282));
    InMux I__9890 (
            .O(N__43299),
            .I(N__43279));
    Span4Mux_v I__9889 (
            .O(N__43296),
            .I(N__43276));
    Span4Mux_v I__9888 (
            .O(N__43293),
            .I(N__43271));
    Span4Mux_h I__9887 (
            .O(N__43290),
            .I(N__43271));
    LocalMux I__9886 (
            .O(N__43287),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    LocalMux I__9885 (
            .O(N__43282),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    LocalMux I__9884 (
            .O(N__43279),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv4 I__9883 (
            .O(N__43276),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv4 I__9882 (
            .O(N__43271),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    CascadeMux I__9881 (
            .O(N__43260),
            .I(N__43254));
    InMux I__9880 (
            .O(N__43259),
            .I(N__43246));
    InMux I__9879 (
            .O(N__43258),
            .I(N__43246));
    InMux I__9878 (
            .O(N__43257),
            .I(N__43243));
    InMux I__9877 (
            .O(N__43254),
            .I(N__43240));
    CascadeMux I__9876 (
            .O(N__43253),
            .I(N__43236));
    InMux I__9875 (
            .O(N__43252),
            .I(N__43229));
    InMux I__9874 (
            .O(N__43251),
            .I(N__43229));
    LocalMux I__9873 (
            .O(N__43246),
            .I(N__43226));
    LocalMux I__9872 (
            .O(N__43243),
            .I(N__43221));
    LocalMux I__9871 (
            .O(N__43240),
            .I(N__43221));
    InMux I__9870 (
            .O(N__43239),
            .I(N__43218));
    InMux I__9869 (
            .O(N__43236),
            .I(N__43215));
    InMux I__9868 (
            .O(N__43235),
            .I(N__43210));
    InMux I__9867 (
            .O(N__43234),
            .I(N__43210));
    LocalMux I__9866 (
            .O(N__43229),
            .I(N__43207));
    Span4Mux_h I__9865 (
            .O(N__43226),
            .I(N__43204));
    Span4Mux_v I__9864 (
            .O(N__43221),
            .I(N__43199));
    LocalMux I__9863 (
            .O(N__43218),
            .I(N__43199));
    LocalMux I__9862 (
            .O(N__43215),
            .I(measured_delay_tr_15));
    LocalMux I__9861 (
            .O(N__43210),
            .I(measured_delay_tr_15));
    Odrv4 I__9860 (
            .O(N__43207),
            .I(measured_delay_tr_15));
    Odrv4 I__9859 (
            .O(N__43204),
            .I(measured_delay_tr_15));
    Odrv4 I__9858 (
            .O(N__43199),
            .I(measured_delay_tr_15));
    CascadeMux I__9857 (
            .O(N__43188),
            .I(N__43185));
    InMux I__9856 (
            .O(N__43185),
            .I(N__43182));
    LocalMux I__9855 (
            .O(N__43182),
            .I(N__43179));
    Span4Mux_h I__9854 (
            .O(N__43179),
            .I(N__43176));
    Odrv4 I__9853 (
            .O(N__43176),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__9852 (
            .O(N__43173),
            .I(N__43170));
    InMux I__9851 (
            .O(N__43170),
            .I(N__43167));
    LocalMux I__9850 (
            .O(N__43167),
            .I(N__43164));
    Span4Mux_h I__9849 (
            .O(N__43164),
            .I(N__43161));
    Odrv4 I__9848 (
            .O(N__43161),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__9847 (
            .O(N__43158),
            .I(N__43149));
    InMux I__9846 (
            .O(N__43157),
            .I(N__43149));
    InMux I__9845 (
            .O(N__43156),
            .I(N__43149));
    LocalMux I__9844 (
            .O(N__43149),
            .I(N__43145));
    InMux I__9843 (
            .O(N__43148),
            .I(N__43142));
    Span4Mux_h I__9842 (
            .O(N__43145),
            .I(N__43134));
    LocalMux I__9841 (
            .O(N__43142),
            .I(N__43131));
    InMux I__9840 (
            .O(N__43141),
            .I(N__43128));
    InMux I__9839 (
            .O(N__43140),
            .I(N__43119));
    InMux I__9838 (
            .O(N__43139),
            .I(N__43119));
    InMux I__9837 (
            .O(N__43138),
            .I(N__43119));
    InMux I__9836 (
            .O(N__43137),
            .I(N__43119));
    Odrv4 I__9835 (
            .O(N__43134),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    Odrv4 I__9834 (
            .O(N__43131),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    LocalMux I__9833 (
            .O(N__43128),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    LocalMux I__9832 (
            .O(N__43119),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    InMux I__9831 (
            .O(N__43110),
            .I(N__43106));
    InMux I__9830 (
            .O(N__43109),
            .I(N__43102));
    LocalMux I__9829 (
            .O(N__43106),
            .I(N__43099));
    InMux I__9828 (
            .O(N__43105),
            .I(N__43096));
    LocalMux I__9827 (
            .O(N__43102),
            .I(N__43093));
    Span4Mux_h I__9826 (
            .O(N__43099),
            .I(N__43088));
    LocalMux I__9825 (
            .O(N__43096),
            .I(N__43088));
    Odrv12 I__9824 (
            .O(N__43093),
            .I(measured_delay_tr_10));
    Odrv4 I__9823 (
            .O(N__43088),
            .I(measured_delay_tr_10));
    CascadeMux I__9822 (
            .O(N__43083),
            .I(N__43080));
    InMux I__9821 (
            .O(N__43080),
            .I(N__43077));
    LocalMux I__9820 (
            .O(N__43077),
            .I(N__43074));
    Span4Mux_v I__9819 (
            .O(N__43074),
            .I(N__43071));
    Odrv4 I__9818 (
            .O(N__43071),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CEMux I__9817 (
            .O(N__43068),
            .I(N__43064));
    CEMux I__9816 (
            .O(N__43067),
            .I(N__43059));
    LocalMux I__9815 (
            .O(N__43064),
            .I(N__43056));
    CEMux I__9814 (
            .O(N__43063),
            .I(N__43053));
    CEMux I__9813 (
            .O(N__43062),
            .I(N__43050));
    LocalMux I__9812 (
            .O(N__43059),
            .I(N__43047));
    Span4Mux_v I__9811 (
            .O(N__43056),
            .I(N__43041));
    LocalMux I__9810 (
            .O(N__43053),
            .I(N__43041));
    LocalMux I__9809 (
            .O(N__43050),
            .I(N__43038));
    Span4Mux_h I__9808 (
            .O(N__43047),
            .I(N__43035));
    CEMux I__9807 (
            .O(N__43046),
            .I(N__43032));
    Span4Mux_v I__9806 (
            .O(N__43041),
            .I(N__43029));
    Span4Mux_v I__9805 (
            .O(N__43038),
            .I(N__43026));
    Span4Mux_v I__9804 (
            .O(N__43035),
            .I(N__43021));
    LocalMux I__9803 (
            .O(N__43032),
            .I(N__43021));
    Span4Mux_h I__9802 (
            .O(N__43029),
            .I(N__43018));
    Span4Mux_h I__9801 (
            .O(N__43026),
            .I(N__43015));
    Span4Mux_h I__9800 (
            .O(N__43021),
            .I(N__43012));
    Odrv4 I__9799 (
            .O(N__43018),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__9798 (
            .O(N__43015),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__9797 (
            .O(N__43012),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__9796 (
            .O(N__43005),
            .I(N__43002));
    LocalMux I__9795 (
            .O(N__43002),
            .I(N__42996));
    InMux I__9794 (
            .O(N__43001),
            .I(N__42993));
    InMux I__9793 (
            .O(N__43000),
            .I(N__42990));
    InMux I__9792 (
            .O(N__42999),
            .I(N__42987));
    Span4Mux_h I__9791 (
            .O(N__42996),
            .I(N__42984));
    LocalMux I__9790 (
            .O(N__42993),
            .I(N__42981));
    LocalMux I__9789 (
            .O(N__42990),
            .I(N__42978));
    LocalMux I__9788 (
            .O(N__42987),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__9787 (
            .O(N__42984),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__9786 (
            .O(N__42981),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__9785 (
            .O(N__42978),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__9784 (
            .O(N__42969),
            .I(N__42964));
    InMux I__9783 (
            .O(N__42968),
            .I(N__42961));
    InMux I__9782 (
            .O(N__42967),
            .I(N__42958));
    LocalMux I__9781 (
            .O(N__42964),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__9780 (
            .O(N__42961),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__9779 (
            .O(N__42958),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__9778 (
            .O(N__42951),
            .I(bfn_18_7_0_));
    InMux I__9777 (
            .O(N__42948),
            .I(N__42943));
    InMux I__9776 (
            .O(N__42947),
            .I(N__42940));
    InMux I__9775 (
            .O(N__42946),
            .I(N__42937));
    LocalMux I__9774 (
            .O(N__42943),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__9773 (
            .O(N__42940),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__9772 (
            .O(N__42937),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__9771 (
            .O(N__42930),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    CascadeMux I__9770 (
            .O(N__42927),
            .I(N__42922));
    InMux I__9769 (
            .O(N__42926),
            .I(N__42919));
    InMux I__9768 (
            .O(N__42925),
            .I(N__42916));
    InMux I__9767 (
            .O(N__42922),
            .I(N__42913));
    LocalMux I__9766 (
            .O(N__42919),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__9765 (
            .O(N__42916),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__9764 (
            .O(N__42913),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__9763 (
            .O(N__42906),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__9762 (
            .O(N__42903),
            .I(N__42898));
    CascadeMux I__9761 (
            .O(N__42902),
            .I(N__42895));
    InMux I__9760 (
            .O(N__42901),
            .I(N__42890));
    LocalMux I__9759 (
            .O(N__42898),
            .I(N__42887));
    InMux I__9758 (
            .O(N__42895),
            .I(N__42884));
    InMux I__9757 (
            .O(N__42894),
            .I(N__42881));
    InMux I__9756 (
            .O(N__42893),
            .I(N__42878));
    LocalMux I__9755 (
            .O(N__42890),
            .I(N__42873));
    Span4Mux_h I__9754 (
            .O(N__42887),
            .I(N__42873));
    LocalMux I__9753 (
            .O(N__42884),
            .I(measured_delay_tr_14));
    LocalMux I__9752 (
            .O(N__42881),
            .I(measured_delay_tr_14));
    LocalMux I__9751 (
            .O(N__42878),
            .I(measured_delay_tr_14));
    Odrv4 I__9750 (
            .O(N__42873),
            .I(measured_delay_tr_14));
    InMux I__9749 (
            .O(N__42864),
            .I(N__42861));
    LocalMux I__9748 (
            .O(N__42861),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ));
    InMux I__9747 (
            .O(N__42858),
            .I(N__42854));
    InMux I__9746 (
            .O(N__42857),
            .I(N__42851));
    LocalMux I__9745 (
            .O(N__42854),
            .I(N__42848));
    LocalMux I__9744 (
            .O(N__42851),
            .I(N__42845));
    Span12Mux_v I__9743 (
            .O(N__42848),
            .I(N__42841));
    Span4Mux_h I__9742 (
            .O(N__42845),
            .I(N__42838));
    InMux I__9741 (
            .O(N__42844),
            .I(N__42835));
    Odrv12 I__9740 (
            .O(N__42841),
            .I(measured_delay_tr_6));
    Odrv4 I__9739 (
            .O(N__42838),
            .I(measured_delay_tr_6));
    LocalMux I__9738 (
            .O(N__42835),
            .I(measured_delay_tr_6));
    CascadeMux I__9737 (
            .O(N__42828),
            .I(N__42825));
    InMux I__9736 (
            .O(N__42825),
            .I(N__42818));
    InMux I__9735 (
            .O(N__42824),
            .I(N__42815));
    InMux I__9734 (
            .O(N__42823),
            .I(N__42808));
    InMux I__9733 (
            .O(N__42822),
            .I(N__42808));
    InMux I__9732 (
            .O(N__42821),
            .I(N__42808));
    LocalMux I__9731 (
            .O(N__42818),
            .I(N__42803));
    LocalMux I__9730 (
            .O(N__42815),
            .I(N__42803));
    LocalMux I__9729 (
            .O(N__42808),
            .I(N__42800));
    Span4Mux_v I__9728 (
            .O(N__42803),
            .I(N__42796));
    Span4Mux_v I__9727 (
            .O(N__42800),
            .I(N__42793));
    InMux I__9726 (
            .O(N__42799),
            .I(N__42790));
    Odrv4 I__9725 (
            .O(N__42796),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ));
    Odrv4 I__9724 (
            .O(N__42793),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ));
    LocalMux I__9723 (
            .O(N__42790),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ));
    CascadeMux I__9722 (
            .O(N__42783),
            .I(N__42778));
    InMux I__9721 (
            .O(N__42782),
            .I(N__42768));
    InMux I__9720 (
            .O(N__42781),
            .I(N__42768));
    InMux I__9719 (
            .O(N__42778),
            .I(N__42761));
    InMux I__9718 (
            .O(N__42777),
            .I(N__42761));
    InMux I__9717 (
            .O(N__42776),
            .I(N__42761));
    InMux I__9716 (
            .O(N__42775),
            .I(N__42758));
    InMux I__9715 (
            .O(N__42774),
            .I(N__42753));
    InMux I__9714 (
            .O(N__42773),
            .I(N__42753));
    LocalMux I__9713 (
            .O(N__42768),
            .I(N__42746));
    LocalMux I__9712 (
            .O(N__42761),
            .I(N__42746));
    LocalMux I__9711 (
            .O(N__42758),
            .I(N__42743));
    LocalMux I__9710 (
            .O(N__42753),
            .I(N__42740));
    InMux I__9709 (
            .O(N__42752),
            .I(N__42736));
    InMux I__9708 (
            .O(N__42751),
            .I(N__42733));
    Span4Mux_h I__9707 (
            .O(N__42746),
            .I(N__42730));
    Span4Mux_v I__9706 (
            .O(N__42743),
            .I(N__42725));
    Span4Mux_v I__9705 (
            .O(N__42740),
            .I(N__42725));
    InMux I__9704 (
            .O(N__42739),
            .I(N__42722));
    LocalMux I__9703 (
            .O(N__42736),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    LocalMux I__9702 (
            .O(N__42733),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    Odrv4 I__9701 (
            .O(N__42730),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    Odrv4 I__9700 (
            .O(N__42725),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    LocalMux I__9699 (
            .O(N__42722),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    CascadeMux I__9698 (
            .O(N__42711),
            .I(N__42708));
    InMux I__9697 (
            .O(N__42708),
            .I(N__42705));
    LocalMux I__9696 (
            .O(N__42705),
            .I(N__42702));
    Odrv4 I__9695 (
            .O(N__42702),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__9694 (
            .O(N__42699),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15_cascade_ ));
    CascadeMux I__9693 (
            .O(N__42696),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_ ));
    CascadeMux I__9692 (
            .O(N__42693),
            .I(N__42690));
    InMux I__9691 (
            .O(N__42690),
            .I(N__42687));
    LocalMux I__9690 (
            .O(N__42687),
            .I(N__42684));
    Odrv4 I__9689 (
            .O(N__42684),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ));
    InMux I__9688 (
            .O(N__42681),
            .I(N__42676));
    InMux I__9687 (
            .O(N__42680),
            .I(N__42673));
    InMux I__9686 (
            .O(N__42679),
            .I(N__42670));
    LocalMux I__9685 (
            .O(N__42676),
            .I(N__42667));
    LocalMux I__9684 (
            .O(N__42673),
            .I(N__42662));
    LocalMux I__9683 (
            .O(N__42670),
            .I(N__42662));
    Odrv12 I__9682 (
            .O(N__42667),
            .I(measured_delay_tr_11));
    Odrv4 I__9681 (
            .O(N__42662),
            .I(measured_delay_tr_11));
    CascadeMux I__9680 (
            .O(N__42657),
            .I(N__42654));
    InMux I__9679 (
            .O(N__42654),
            .I(N__42651));
    LocalMux I__9678 (
            .O(N__42651),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ));
    InMux I__9677 (
            .O(N__42648),
            .I(N__42643));
    InMux I__9676 (
            .O(N__42647),
            .I(N__42640));
    InMux I__9675 (
            .O(N__42646),
            .I(N__42637));
    LocalMux I__9674 (
            .O(N__42643),
            .I(N__42634));
    LocalMux I__9673 (
            .O(N__42640),
            .I(N__42629));
    LocalMux I__9672 (
            .O(N__42637),
            .I(N__42629));
    Odrv12 I__9671 (
            .O(N__42634),
            .I(measured_delay_tr_12));
    Odrv4 I__9670 (
            .O(N__42629),
            .I(measured_delay_tr_12));
    CascadeMux I__9669 (
            .O(N__42624),
            .I(N__42621));
    InMux I__9668 (
            .O(N__42621),
            .I(N__42618));
    LocalMux I__9667 (
            .O(N__42618),
            .I(N__42615));
    Odrv12 I__9666 (
            .O(N__42615),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__9665 (
            .O(N__42612),
            .I(N__42608));
    InMux I__9664 (
            .O(N__42611),
            .I(N__42604));
    InMux I__9663 (
            .O(N__42608),
            .I(N__42601));
    InMux I__9662 (
            .O(N__42607),
            .I(N__42598));
    LocalMux I__9661 (
            .O(N__42604),
            .I(N__42595));
    LocalMux I__9660 (
            .O(N__42601),
            .I(N__42592));
    LocalMux I__9659 (
            .O(N__42598),
            .I(N__42589));
    Span4Mux_v I__9658 (
            .O(N__42595),
            .I(N__42584));
    Span4Mux_h I__9657 (
            .O(N__42592),
            .I(N__42584));
    Odrv12 I__9656 (
            .O(N__42589),
            .I(measured_delay_tr_13));
    Odrv4 I__9655 (
            .O(N__42584),
            .I(measured_delay_tr_13));
    CascadeMux I__9654 (
            .O(N__42579),
            .I(N__42576));
    InMux I__9653 (
            .O(N__42576),
            .I(N__42573));
    LocalMux I__9652 (
            .O(N__42573),
            .I(N__42570));
    Odrv4 I__9651 (
            .O(N__42570),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ));
    InMux I__9650 (
            .O(N__42567),
            .I(N__42564));
    LocalMux I__9649 (
            .O(N__42564),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    InMux I__9648 (
            .O(N__42561),
            .I(N__42558));
    LocalMux I__9647 (
            .O(N__42558),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__9646 (
            .O(N__42555),
            .I(N__42552));
    LocalMux I__9645 (
            .O(N__42552),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__9644 (
            .O(N__42549),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__9643 (
            .O(N__42546),
            .I(N__42543));
    InMux I__9642 (
            .O(N__42543),
            .I(N__42540));
    LocalMux I__9641 (
            .O(N__42540),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__9640 (
            .O(N__42537),
            .I(N__42534));
    InMux I__9639 (
            .O(N__42534),
            .I(N__42531));
    LocalMux I__9638 (
            .O(N__42531),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__9637 (
            .O(N__42528),
            .I(N__42525));
    InMux I__9636 (
            .O(N__42525),
            .I(N__42522));
    LocalMux I__9635 (
            .O(N__42522),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__9634 (
            .O(N__42519),
            .I(N__42516));
    InMux I__9633 (
            .O(N__42516),
            .I(N__42513));
    LocalMux I__9632 (
            .O(N__42513),
            .I(N__42510));
    Odrv4 I__9631 (
            .O(N__42510),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ));
    InMux I__9630 (
            .O(N__42507),
            .I(N__42503));
    InMux I__9629 (
            .O(N__42506),
            .I(N__42500));
    LocalMux I__9628 (
            .O(N__42503),
            .I(N__42497));
    LocalMux I__9627 (
            .O(N__42500),
            .I(N__42494));
    Span4Mux_h I__9626 (
            .O(N__42497),
            .I(N__42490));
    Span4Mux_h I__9625 (
            .O(N__42494),
            .I(N__42487));
    InMux I__9624 (
            .O(N__42493),
            .I(N__42484));
    Odrv4 I__9623 (
            .O(N__42490),
            .I(measured_delay_tr_7));
    Odrv4 I__9622 (
            .O(N__42487),
            .I(measured_delay_tr_7));
    LocalMux I__9621 (
            .O(N__42484),
            .I(measured_delay_tr_7));
    CascadeMux I__9620 (
            .O(N__42477),
            .I(N__42474));
    InMux I__9619 (
            .O(N__42474),
            .I(N__42471));
    LocalMux I__9618 (
            .O(N__42471),
            .I(N__42468));
    Odrv4 I__9617 (
            .O(N__42468),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__9616 (
            .O(N__42465),
            .I(N__42462));
    InMux I__9615 (
            .O(N__42462),
            .I(N__42459));
    LocalMux I__9614 (
            .O(N__42459),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__9613 (
            .O(N__42456),
            .I(N__42453));
    LocalMux I__9612 (
            .O(N__42453),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__9611 (
            .O(N__42450),
            .I(N__42447));
    LocalMux I__9610 (
            .O(N__42447),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__9609 (
            .O(N__42444),
            .I(N__42441));
    InMux I__9608 (
            .O(N__42441),
            .I(N__42438));
    LocalMux I__9607 (
            .O(N__42438),
            .I(N__42435));
    Odrv12 I__9606 (
            .O(N__42435),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__9605 (
            .O(N__42432),
            .I(N__42429));
    LocalMux I__9604 (
            .O(N__42429),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__9603 (
            .O(N__42426),
            .I(N__42423));
    InMux I__9602 (
            .O(N__42423),
            .I(N__42420));
    LocalMux I__9601 (
            .O(N__42420),
            .I(N__42417));
    Odrv12 I__9600 (
            .O(N__42417),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    InMux I__9599 (
            .O(N__42414),
            .I(N__42411));
    LocalMux I__9598 (
            .O(N__42411),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__9597 (
            .O(N__42408),
            .I(N__42405));
    InMux I__9596 (
            .O(N__42405),
            .I(N__42402));
    LocalMux I__9595 (
            .O(N__42402),
            .I(N__42399));
    Span4Mux_h I__9594 (
            .O(N__42399),
            .I(N__42396));
    Odrv4 I__9593 (
            .O(N__42396),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__9592 (
            .O(N__42393),
            .I(N__42390));
    LocalMux I__9591 (
            .O(N__42390),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__9590 (
            .O(N__42387),
            .I(N__42384));
    InMux I__9589 (
            .O(N__42384),
            .I(N__42381));
    LocalMux I__9588 (
            .O(N__42381),
            .I(N__42378));
    Odrv4 I__9587 (
            .O(N__42378),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__9586 (
            .O(N__42375),
            .I(N__42372));
    LocalMux I__9585 (
            .O(N__42372),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__9584 (
            .O(N__42369),
            .I(N__42366));
    LocalMux I__9583 (
            .O(N__42366),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__9582 (
            .O(N__42363),
            .I(N__42360));
    LocalMux I__9581 (
            .O(N__42360),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__9580 (
            .O(N__42357),
            .I(N__42354));
    InMux I__9579 (
            .O(N__42354),
            .I(N__42351));
    LocalMux I__9578 (
            .O(N__42351),
            .I(N__42348));
    Odrv4 I__9577 (
            .O(N__42348),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__9576 (
            .O(N__42345),
            .I(N__42342));
    LocalMux I__9575 (
            .O(N__42342),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__9574 (
            .O(N__42339),
            .I(N__42336));
    InMux I__9573 (
            .O(N__42336),
            .I(N__42333));
    LocalMux I__9572 (
            .O(N__42333),
            .I(N__42330));
    Span4Mux_v I__9571 (
            .O(N__42330),
            .I(N__42327));
    Odrv4 I__9570 (
            .O(N__42327),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    InMux I__9569 (
            .O(N__42324),
            .I(N__42321));
    LocalMux I__9568 (
            .O(N__42321),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__9567 (
            .O(N__42318),
            .I(N__42315));
    InMux I__9566 (
            .O(N__42315),
            .I(N__42312));
    LocalMux I__9565 (
            .O(N__42312),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__9564 (
            .O(N__42309),
            .I(N__42306));
    LocalMux I__9563 (
            .O(N__42306),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__9562 (
            .O(N__42303),
            .I(N__42300));
    InMux I__9561 (
            .O(N__42300),
            .I(N__42297));
    LocalMux I__9560 (
            .O(N__42297),
            .I(N__42294));
    Odrv4 I__9559 (
            .O(N__42294),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__9558 (
            .O(N__42291),
            .I(N__42288));
    LocalMux I__9557 (
            .O(N__42288),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__9556 (
            .O(N__42285),
            .I(N__42282));
    InMux I__9555 (
            .O(N__42282),
            .I(N__42279));
    LocalMux I__9554 (
            .O(N__42279),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__9553 (
            .O(N__42276),
            .I(N__42273));
    LocalMux I__9552 (
            .O(N__42273),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__9551 (
            .O(N__42270),
            .I(N__42267));
    InMux I__9550 (
            .O(N__42267),
            .I(N__42264));
    LocalMux I__9549 (
            .O(N__42264),
            .I(N__42261));
    Odrv4 I__9548 (
            .O(N__42261),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__9547 (
            .O(N__42258),
            .I(N__42255));
    LocalMux I__9546 (
            .O(N__42255),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__9545 (
            .O(N__42252),
            .I(N__42249));
    LocalMux I__9544 (
            .O(N__42249),
            .I(N__42246));
    Span4Mux_h I__9543 (
            .O(N__42246),
            .I(N__42243));
    Odrv4 I__9542 (
            .O(N__42243),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__9541 (
            .O(N__42240),
            .I(N__42237));
    InMux I__9540 (
            .O(N__42237),
            .I(N__42234));
    LocalMux I__9539 (
            .O(N__42234),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__9538 (
            .O(N__42231),
            .I(N__42227));
    CascadeMux I__9537 (
            .O(N__42230),
            .I(N__42214));
    InMux I__9536 (
            .O(N__42227),
            .I(N__42209));
    InMux I__9535 (
            .O(N__42226),
            .I(N__42209));
    CascadeMux I__9534 (
            .O(N__42225),
            .I(N__42202));
    CascadeMux I__9533 (
            .O(N__42224),
            .I(N__42199));
    CascadeMux I__9532 (
            .O(N__42223),
            .I(N__42196));
    CascadeMux I__9531 (
            .O(N__42222),
            .I(N__42193));
    CascadeMux I__9530 (
            .O(N__42221),
            .I(N__42189));
    CascadeMux I__9529 (
            .O(N__42220),
            .I(N__42186));
    CascadeMux I__9528 (
            .O(N__42219),
            .I(N__42183));
    CascadeMux I__9527 (
            .O(N__42218),
            .I(N__42180));
    InMux I__9526 (
            .O(N__42217),
            .I(N__42171));
    InMux I__9525 (
            .O(N__42214),
            .I(N__42171));
    LocalMux I__9524 (
            .O(N__42209),
            .I(N__42168));
    InMux I__9523 (
            .O(N__42208),
            .I(N__42151));
    InMux I__9522 (
            .O(N__42207),
            .I(N__42151));
    InMux I__9521 (
            .O(N__42206),
            .I(N__42151));
    InMux I__9520 (
            .O(N__42205),
            .I(N__42151));
    InMux I__9519 (
            .O(N__42202),
            .I(N__42151));
    InMux I__9518 (
            .O(N__42199),
            .I(N__42151));
    InMux I__9517 (
            .O(N__42196),
            .I(N__42151));
    InMux I__9516 (
            .O(N__42193),
            .I(N__42151));
    CascadeMux I__9515 (
            .O(N__42192),
            .I(N__42148));
    InMux I__9514 (
            .O(N__42189),
            .I(N__42131));
    InMux I__9513 (
            .O(N__42186),
            .I(N__42131));
    InMux I__9512 (
            .O(N__42183),
            .I(N__42131));
    InMux I__9511 (
            .O(N__42180),
            .I(N__42131));
    InMux I__9510 (
            .O(N__42179),
            .I(N__42131));
    InMux I__9509 (
            .O(N__42178),
            .I(N__42131));
    InMux I__9508 (
            .O(N__42177),
            .I(N__42131));
    InMux I__9507 (
            .O(N__42176),
            .I(N__42131));
    LocalMux I__9506 (
            .O(N__42171),
            .I(N__42122));
    Span4Mux_v I__9505 (
            .O(N__42168),
            .I(N__42122));
    LocalMux I__9504 (
            .O(N__42151),
            .I(N__42122));
    InMux I__9503 (
            .O(N__42148),
            .I(N__42119));
    LocalMux I__9502 (
            .O(N__42131),
            .I(N__42116));
    InMux I__9501 (
            .O(N__42130),
            .I(N__42112));
    InMux I__9500 (
            .O(N__42129),
            .I(N__42109));
    Span4Mux_h I__9499 (
            .O(N__42122),
            .I(N__42106));
    LocalMux I__9498 (
            .O(N__42119),
            .I(N__42101));
    Span4Mux_v I__9497 (
            .O(N__42116),
            .I(N__42101));
    InMux I__9496 (
            .O(N__42115),
            .I(N__42098));
    LocalMux I__9495 (
            .O(N__42112),
            .I(N__42095));
    LocalMux I__9494 (
            .O(N__42109),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9493 (
            .O(N__42106),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9492 (
            .O(N__42101),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    LocalMux I__9491 (
            .O(N__42098),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv12 I__9490 (
            .O(N__42095),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    InMux I__9489 (
            .O(N__42084),
            .I(N__42081));
    LocalMux I__9488 (
            .O(N__42081),
            .I(N__42078));
    Span4Mux_h I__9487 (
            .O(N__42078),
            .I(N__42075));
    Odrv4 I__9486 (
            .O(N__42075),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    InMux I__9485 (
            .O(N__42072),
            .I(N__42068));
    InMux I__9484 (
            .O(N__42071),
            .I(N__42065));
    LocalMux I__9483 (
            .O(N__42068),
            .I(N__42062));
    LocalMux I__9482 (
            .O(N__42065),
            .I(N__42059));
    Span4Mux_h I__9481 (
            .O(N__42062),
            .I(N__42056));
    Span4Mux_v I__9480 (
            .O(N__42059),
            .I(N__42051));
    Span4Mux_v I__9479 (
            .O(N__42056),
            .I(N__42048));
    InMux I__9478 (
            .O(N__42055),
            .I(N__42045));
    InMux I__9477 (
            .O(N__42054),
            .I(N__42042));
    Odrv4 I__9476 (
            .O(N__42051),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    Odrv4 I__9475 (
            .O(N__42048),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__9474 (
            .O(N__42045),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__9473 (
            .O(N__42042),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    InMux I__9472 (
            .O(N__42033),
            .I(N__42030));
    LocalMux I__9471 (
            .O(N__42030),
            .I(N__42026));
    InMux I__9470 (
            .O(N__42029),
            .I(N__42023));
    Span4Mux_h I__9469 (
            .O(N__42026),
            .I(N__42020));
    LocalMux I__9468 (
            .O(N__42023),
            .I(N__42017));
    Odrv4 I__9467 (
            .O(N__42020),
            .I(\phase_controller_inst1.N_231 ));
    Odrv4 I__9466 (
            .O(N__42017),
            .I(\phase_controller_inst1.N_231 ));
    CascadeMux I__9465 (
            .O(N__42012),
            .I(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_ ));
    InMux I__9464 (
            .O(N__42009),
            .I(N__42004));
    InMux I__9463 (
            .O(N__42008),
            .I(N__42001));
    InMux I__9462 (
            .O(N__42007),
            .I(N__41998));
    LocalMux I__9461 (
            .O(N__42004),
            .I(N__41990));
    LocalMux I__9460 (
            .O(N__42001),
            .I(N__41990));
    LocalMux I__9459 (
            .O(N__41998),
            .I(N__41990));
    InMux I__9458 (
            .O(N__41997),
            .I(N__41987));
    Span4Mux_v I__9457 (
            .O(N__41990),
            .I(N__41984));
    LocalMux I__9456 (
            .O(N__41987),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv4 I__9455 (
            .O(N__41984),
            .I(\phase_controller_inst1.tr_time_passed ));
    CascadeMux I__9454 (
            .O(N__41979),
            .I(N__41976));
    InMux I__9453 (
            .O(N__41976),
            .I(N__41973));
    LocalMux I__9452 (
            .O(N__41973),
            .I(N__41970));
    Odrv4 I__9451 (
            .O(N__41970),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__9450 (
            .O(N__41967),
            .I(N__41964));
    LocalMux I__9449 (
            .O(N__41964),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__9448 (
            .O(N__41961),
            .I(N__41958));
    LocalMux I__9447 (
            .O(N__41958),
            .I(N__41954));
    InMux I__9446 (
            .O(N__41957),
            .I(N__41951));
    Odrv12 I__9445 (
            .O(N__41954),
            .I(\delay_measurement_inst.elapsed_time_hc_26 ));
    LocalMux I__9444 (
            .O(N__41951),
            .I(\delay_measurement_inst.elapsed_time_hc_26 ));
    InMux I__9443 (
            .O(N__41946),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__9442 (
            .O(N__41943),
            .I(N__41940));
    LocalMux I__9441 (
            .O(N__41940),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__9440 (
            .O(N__41937),
            .I(bfn_17_11_0_));
    InMux I__9439 (
            .O(N__41934),
            .I(N__41931));
    LocalMux I__9438 (
            .O(N__41931),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__9437 (
            .O(N__41928),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__9436 (
            .O(N__41925),
            .I(N__41922));
    LocalMux I__9435 (
            .O(N__41922),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__9434 (
            .O(N__41919),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__9433 (
            .O(N__41916),
            .I(N__41913));
    InMux I__9432 (
            .O(N__41913),
            .I(N__41910));
    LocalMux I__9431 (
            .O(N__41910),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ));
    InMux I__9430 (
            .O(N__41907),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__9429 (
            .O(N__41904),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__9428 (
            .O(N__41901),
            .I(N__41896));
    CascadeMux I__9427 (
            .O(N__41900),
            .I(N__41889));
    CascadeMux I__9426 (
            .O(N__41899),
            .I(N__41886));
    InMux I__9425 (
            .O(N__41896),
            .I(N__41881));
    InMux I__9424 (
            .O(N__41895),
            .I(N__41881));
    CascadeMux I__9423 (
            .O(N__41894),
            .I(N__41876));
    CascadeMux I__9422 (
            .O(N__41893),
            .I(N__41873));
    CascadeMux I__9421 (
            .O(N__41892),
            .I(N__41870));
    InMux I__9420 (
            .O(N__41889),
            .I(N__41866));
    InMux I__9419 (
            .O(N__41886),
            .I(N__41863));
    LocalMux I__9418 (
            .O(N__41881),
            .I(N__41860));
    InMux I__9417 (
            .O(N__41880),
            .I(N__41857));
    InMux I__9416 (
            .O(N__41879),
            .I(N__41854));
    InMux I__9415 (
            .O(N__41876),
            .I(N__41849));
    InMux I__9414 (
            .O(N__41873),
            .I(N__41842));
    InMux I__9413 (
            .O(N__41870),
            .I(N__41842));
    InMux I__9412 (
            .O(N__41869),
            .I(N__41842));
    LocalMux I__9411 (
            .O(N__41866),
            .I(N__41839));
    LocalMux I__9410 (
            .O(N__41863),
            .I(N__41836));
    Span4Mux_v I__9409 (
            .O(N__41860),
            .I(N__41831));
    LocalMux I__9408 (
            .O(N__41857),
            .I(N__41831));
    LocalMux I__9407 (
            .O(N__41854),
            .I(N__41828));
    InMux I__9406 (
            .O(N__41853),
            .I(N__41825));
    CascadeMux I__9405 (
            .O(N__41852),
            .I(N__41821));
    LocalMux I__9404 (
            .O(N__41849),
            .I(N__41818));
    LocalMux I__9403 (
            .O(N__41842),
            .I(N__41815));
    Span4Mux_v I__9402 (
            .O(N__41839),
            .I(N__41812));
    Span4Mux_h I__9401 (
            .O(N__41836),
            .I(N__41807));
    Span4Mux_h I__9400 (
            .O(N__41831),
            .I(N__41807));
    Span4Mux_v I__9399 (
            .O(N__41828),
            .I(N__41802));
    LocalMux I__9398 (
            .O(N__41825),
            .I(N__41802));
    InMux I__9397 (
            .O(N__41824),
            .I(N__41799));
    InMux I__9396 (
            .O(N__41821),
            .I(N__41795));
    Span4Mux_v I__9395 (
            .O(N__41818),
            .I(N__41790));
    Span4Mux_v I__9394 (
            .O(N__41815),
            .I(N__41790));
    Span4Mux_h I__9393 (
            .O(N__41812),
            .I(N__41785));
    Span4Mux_v I__9392 (
            .O(N__41807),
            .I(N__41785));
    Span4Mux_v I__9391 (
            .O(N__41802),
            .I(N__41780));
    LocalMux I__9390 (
            .O(N__41799),
            .I(N__41780));
    CascadeMux I__9389 (
            .O(N__41798),
            .I(N__41777));
    LocalMux I__9388 (
            .O(N__41795),
            .I(N__41774));
    Span4Mux_h I__9387 (
            .O(N__41790),
            .I(N__41771));
    Span4Mux_h I__9386 (
            .O(N__41785),
            .I(N__41768));
    Span4Mux_h I__9385 (
            .O(N__41780),
            .I(N__41765));
    InMux I__9384 (
            .O(N__41777),
            .I(N__41762));
    Odrv12 I__9383 (
            .O(N__41774),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    Odrv4 I__9382 (
            .O(N__41771),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    Odrv4 I__9381 (
            .O(N__41768),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    Odrv4 I__9380 (
            .O(N__41765),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    LocalMux I__9379 (
            .O(N__41762),
            .I(\delay_measurement_inst.elapsed_time_hc_31 ));
    CEMux I__9378 (
            .O(N__41751),
            .I(N__41736));
    CEMux I__9377 (
            .O(N__41750),
            .I(N__41736));
    CEMux I__9376 (
            .O(N__41749),
            .I(N__41736));
    CEMux I__9375 (
            .O(N__41748),
            .I(N__41736));
    CEMux I__9374 (
            .O(N__41747),
            .I(N__41736));
    GlobalMux I__9373 (
            .O(N__41736),
            .I(N__41733));
    gio2CtrlBuf I__9372 (
            .O(N__41733),
            .I(\delay_measurement_inst.delay_hc_timer.N_335_i_g ));
    InMux I__9371 (
            .O(N__41730),
            .I(N__41727));
    LocalMux I__9370 (
            .O(N__41727),
            .I(N__41722));
    InMux I__9369 (
            .O(N__41726),
            .I(N__41717));
    InMux I__9368 (
            .O(N__41725),
            .I(N__41717));
    Odrv4 I__9367 (
            .O(N__41722),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__9366 (
            .O(N__41717),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    InMux I__9365 (
            .O(N__41712),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__9364 (
            .O(N__41709),
            .I(N__41706));
    LocalMux I__9363 (
            .O(N__41706),
            .I(N__41701));
    InMux I__9362 (
            .O(N__41705),
            .I(N__41698));
    CascadeMux I__9361 (
            .O(N__41704),
            .I(N__41695));
    Span4Mux_h I__9360 (
            .O(N__41701),
            .I(N__41692));
    LocalMux I__9359 (
            .O(N__41698),
            .I(N__41689));
    InMux I__9358 (
            .O(N__41695),
            .I(N__41686));
    Odrv4 I__9357 (
            .O(N__41692),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    Odrv4 I__9356 (
            .O(N__41689),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    LocalMux I__9355 (
            .O(N__41686),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    InMux I__9354 (
            .O(N__41679),
            .I(bfn_17_10_0_));
    InMux I__9353 (
            .O(N__41676),
            .I(N__41670));
    InMux I__9352 (
            .O(N__41675),
            .I(N__41670));
    LocalMux I__9351 (
            .O(N__41670),
            .I(N__41667));
    Odrv4 I__9350 (
            .O(N__41667),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__9349 (
            .O(N__41664),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__9348 (
            .O(N__41661),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__9347 (
            .O(N__41658),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__9346 (
            .O(N__41655),
            .I(N__41652));
    LocalMux I__9345 (
            .O(N__41652),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__9344 (
            .O(N__41649),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__9343 (
            .O(N__41646),
            .I(N__41643));
    LocalMux I__9342 (
            .O(N__41643),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_24 ));
    InMux I__9341 (
            .O(N__41640),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__9340 (
            .O(N__41637),
            .I(N__41634));
    LocalMux I__9339 (
            .O(N__41634),
            .I(N__41631));
    Span4Mux_h I__9338 (
            .O(N__41631),
            .I(N__41627));
    InMux I__9337 (
            .O(N__41630),
            .I(N__41624));
    Odrv4 I__9336 (
            .O(N__41627),
            .I(\delay_measurement_inst.elapsed_time_hc_25 ));
    LocalMux I__9335 (
            .O(N__41624),
            .I(\delay_measurement_inst.elapsed_time_hc_25 ));
    InMux I__9334 (
            .O(N__41619),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__9333 (
            .O(N__41616),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__9332 (
            .O(N__41613),
            .I(N__41610));
    LocalMux I__9331 (
            .O(N__41610),
            .I(N__41606));
    CascadeMux I__9330 (
            .O(N__41609),
            .I(N__41603));
    Span4Mux_h I__9329 (
            .O(N__41606),
            .I(N__41599));
    InMux I__9328 (
            .O(N__41603),
            .I(N__41596));
    InMux I__9327 (
            .O(N__41602),
            .I(N__41593));
    Odrv4 I__9326 (
            .O(N__41599),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    LocalMux I__9325 (
            .O(N__41596),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    LocalMux I__9324 (
            .O(N__41593),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__9323 (
            .O(N__41586),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__9322 (
            .O(N__41583),
            .I(N__41580));
    LocalMux I__9321 (
            .O(N__41580),
            .I(N__41576));
    InMux I__9320 (
            .O(N__41579),
            .I(N__41573));
    Span4Mux_h I__9319 (
            .O(N__41576),
            .I(N__41569));
    LocalMux I__9318 (
            .O(N__41573),
            .I(N__41566));
    InMux I__9317 (
            .O(N__41572),
            .I(N__41563));
    Odrv4 I__9316 (
            .O(N__41569),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    Odrv4 I__9315 (
            .O(N__41566),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    LocalMux I__9314 (
            .O(N__41563),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__9313 (
            .O(N__41556),
            .I(bfn_17_9_0_));
    InMux I__9312 (
            .O(N__41553),
            .I(N__41550));
    LocalMux I__9311 (
            .O(N__41550),
            .I(N__41546));
    CascadeMux I__9310 (
            .O(N__41549),
            .I(N__41543));
    Span4Mux_h I__9309 (
            .O(N__41546),
            .I(N__41539));
    InMux I__9308 (
            .O(N__41543),
            .I(N__41536));
    InMux I__9307 (
            .O(N__41542),
            .I(N__41533));
    Odrv4 I__9306 (
            .O(N__41539),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    LocalMux I__9305 (
            .O(N__41536),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    LocalMux I__9304 (
            .O(N__41533),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    InMux I__9303 (
            .O(N__41526),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__9302 (
            .O(N__41523),
            .I(N__41519));
    CascadeMux I__9301 (
            .O(N__41522),
            .I(N__41515));
    LocalMux I__9300 (
            .O(N__41519),
            .I(N__41512));
    InMux I__9299 (
            .O(N__41518),
            .I(N__41509));
    InMux I__9298 (
            .O(N__41515),
            .I(N__41506));
    Odrv4 I__9297 (
            .O(N__41512),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    LocalMux I__9296 (
            .O(N__41509),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    LocalMux I__9295 (
            .O(N__41506),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    InMux I__9294 (
            .O(N__41499),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__9293 (
            .O(N__41496),
            .I(N__41493));
    LocalMux I__9292 (
            .O(N__41493),
            .I(N__41487));
    InMux I__9291 (
            .O(N__41492),
            .I(N__41482));
    InMux I__9290 (
            .O(N__41491),
            .I(N__41482));
    InMux I__9289 (
            .O(N__41490),
            .I(N__41479));
    Odrv4 I__9288 (
            .O(N__41487),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__9287 (
            .O(N__41482),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__9286 (
            .O(N__41479),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    InMux I__9285 (
            .O(N__41472),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__9284 (
            .O(N__41469),
            .I(N__41466));
    LocalMux I__9283 (
            .O(N__41466),
            .I(N__41457));
    InMux I__9282 (
            .O(N__41465),
            .I(N__41450));
    InMux I__9281 (
            .O(N__41464),
            .I(N__41450));
    InMux I__9280 (
            .O(N__41463),
            .I(N__41450));
    InMux I__9279 (
            .O(N__41462),
            .I(N__41443));
    InMux I__9278 (
            .O(N__41461),
            .I(N__41443));
    InMux I__9277 (
            .O(N__41460),
            .I(N__41443));
    Odrv4 I__9276 (
            .O(N__41457),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__9275 (
            .O(N__41450),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__9274 (
            .O(N__41443),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    InMux I__9273 (
            .O(N__41436),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__9272 (
            .O(N__41433),
            .I(N__41430));
    LocalMux I__9271 (
            .O(N__41430),
            .I(N__41425));
    InMux I__9270 (
            .O(N__41429),
            .I(N__41422));
    InMux I__9269 (
            .O(N__41428),
            .I(N__41419));
    Odrv4 I__9268 (
            .O(N__41425),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    LocalMux I__9267 (
            .O(N__41422),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    LocalMux I__9266 (
            .O(N__41419),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    InMux I__9265 (
            .O(N__41412),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__9264 (
            .O(N__41409),
            .I(N__41406));
    LocalMux I__9263 (
            .O(N__41406),
            .I(N__41401));
    InMux I__9262 (
            .O(N__41405),
            .I(N__41396));
    InMux I__9261 (
            .O(N__41404),
            .I(N__41396));
    Odrv4 I__9260 (
            .O(N__41401),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    LocalMux I__9259 (
            .O(N__41396),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    InMux I__9258 (
            .O(N__41391),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__9257 (
            .O(N__41388),
            .I(N__41385));
    InMux I__9256 (
            .O(N__41385),
            .I(N__41382));
    LocalMux I__9255 (
            .O(N__41382),
            .I(N__41379));
    Span4Mux_v I__9254 (
            .O(N__41379),
            .I(N__41375));
    InMux I__9253 (
            .O(N__41378),
            .I(N__41372));
    Odrv4 I__9252 (
            .O(N__41375),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    LocalMux I__9251 (
            .O(N__41372),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    CascadeMux I__9250 (
            .O(N__41367),
            .I(N__41364));
    InMux I__9249 (
            .O(N__41364),
            .I(N__41359));
    InMux I__9248 (
            .O(N__41363),
            .I(N__41356));
    InMux I__9247 (
            .O(N__41362),
            .I(N__41353));
    LocalMux I__9246 (
            .O(N__41359),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    LocalMux I__9245 (
            .O(N__41356),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    LocalMux I__9244 (
            .O(N__41353),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    CascadeMux I__9243 (
            .O(N__41346),
            .I(N__41343));
    InMux I__9242 (
            .O(N__41343),
            .I(N__41340));
    LocalMux I__9241 (
            .O(N__41340),
            .I(N__41337));
    Span4Mux_h I__9240 (
            .O(N__41337),
            .I(N__41332));
    InMux I__9239 (
            .O(N__41336),
            .I(N__41329));
    InMux I__9238 (
            .O(N__41335),
            .I(N__41326));
    Odrv4 I__9237 (
            .O(N__41332),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__9236 (
            .O(N__41329),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__9235 (
            .O(N__41326),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    CascadeMux I__9234 (
            .O(N__41319),
            .I(N__41316));
    InMux I__9233 (
            .O(N__41316),
            .I(N__41313));
    LocalMux I__9232 (
            .O(N__41313),
            .I(N__41309));
    CascadeMux I__9231 (
            .O(N__41312),
            .I(N__41306));
    Span4Mux_h I__9230 (
            .O(N__41309),
            .I(N__41302));
    InMux I__9229 (
            .O(N__41306),
            .I(N__41297));
    InMux I__9228 (
            .O(N__41305),
            .I(N__41297));
    Odrv4 I__9227 (
            .O(N__41302),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    LocalMux I__9226 (
            .O(N__41297),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    InMux I__9225 (
            .O(N__41292),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__9224 (
            .O(N__41289),
            .I(N__41286));
    LocalMux I__9223 (
            .O(N__41286),
            .I(N__41282));
    CascadeMux I__9222 (
            .O(N__41285),
            .I(N__41278));
    Span4Mux_h I__9221 (
            .O(N__41282),
            .I(N__41275));
    InMux I__9220 (
            .O(N__41281),
            .I(N__41272));
    InMux I__9219 (
            .O(N__41278),
            .I(N__41269));
    Odrv4 I__9218 (
            .O(N__41275),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    LocalMux I__9217 (
            .O(N__41272),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    LocalMux I__9216 (
            .O(N__41269),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    InMux I__9215 (
            .O(N__41262),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__9214 (
            .O(N__41259),
            .I(N__41254));
    CascadeMux I__9213 (
            .O(N__41258),
            .I(N__41251));
    CascadeMux I__9212 (
            .O(N__41257),
            .I(N__41247));
    LocalMux I__9211 (
            .O(N__41254),
            .I(N__41244));
    InMux I__9210 (
            .O(N__41251),
            .I(N__41239));
    InMux I__9209 (
            .O(N__41250),
            .I(N__41239));
    InMux I__9208 (
            .O(N__41247),
            .I(N__41236));
    Span4Mux_h I__9207 (
            .O(N__41244),
            .I(N__41233));
    LocalMux I__9206 (
            .O(N__41239),
            .I(N__41228));
    LocalMux I__9205 (
            .O(N__41236),
            .I(N__41228));
    Odrv4 I__9204 (
            .O(N__41233),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    Odrv4 I__9203 (
            .O(N__41228),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    InMux I__9202 (
            .O(N__41223),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__9201 (
            .O(N__41220),
            .I(N__41217));
    LocalMux I__9200 (
            .O(N__41217),
            .I(N__41214));
    Span4Mux_h I__9199 (
            .O(N__41214),
            .I(N__41207));
    InMux I__9198 (
            .O(N__41213),
            .I(N__41200));
    InMux I__9197 (
            .O(N__41212),
            .I(N__41200));
    InMux I__9196 (
            .O(N__41211),
            .I(N__41200));
    InMux I__9195 (
            .O(N__41210),
            .I(N__41197));
    Odrv4 I__9194 (
            .O(N__41207),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__9193 (
            .O(N__41200),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__9192 (
            .O(N__41197),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    InMux I__9191 (
            .O(N__41190),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__9190 (
            .O(N__41187),
            .I(N__41183));
    CascadeMux I__9189 (
            .O(N__41186),
            .I(N__41177));
    LocalMux I__9188 (
            .O(N__41183),
            .I(N__41174));
    InMux I__9187 (
            .O(N__41182),
            .I(N__41167));
    InMux I__9186 (
            .O(N__41181),
            .I(N__41167));
    InMux I__9185 (
            .O(N__41180),
            .I(N__41167));
    InMux I__9184 (
            .O(N__41177),
            .I(N__41164));
    Odrv4 I__9183 (
            .O(N__41174),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__9182 (
            .O(N__41167),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__9181 (
            .O(N__41164),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    InMux I__9180 (
            .O(N__41157),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__9179 (
            .O(N__41154),
            .I(N__41151));
    LocalMux I__9178 (
            .O(N__41151),
            .I(N__41146));
    CascadeMux I__9177 (
            .O(N__41150),
            .I(N__41142));
    CascadeMux I__9176 (
            .O(N__41149),
            .I(N__41139));
    Span4Mux_h I__9175 (
            .O(N__41146),
            .I(N__41136));
    InMux I__9174 (
            .O(N__41145),
            .I(N__41133));
    InMux I__9173 (
            .O(N__41142),
            .I(N__41130));
    InMux I__9172 (
            .O(N__41139),
            .I(N__41127));
    Odrv4 I__9171 (
            .O(N__41136),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__9170 (
            .O(N__41133),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__9169 (
            .O(N__41130),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__9168 (
            .O(N__41127),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    InMux I__9167 (
            .O(N__41118),
            .I(N__41115));
    LocalMux I__9166 (
            .O(N__41115),
            .I(N__41111));
    InMux I__9165 (
            .O(N__41114),
            .I(N__41108));
    Span4Mux_v I__9164 (
            .O(N__41111),
            .I(N__41105));
    LocalMux I__9163 (
            .O(N__41108),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__9162 (
            .O(N__41105),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__9161 (
            .O(N__41100),
            .I(N__41097));
    LocalMux I__9160 (
            .O(N__41097),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ));
    InMux I__9159 (
            .O(N__41094),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__9158 (
            .O(N__41091),
            .I(N__41086));
    InMux I__9157 (
            .O(N__41090),
            .I(N__41081));
    InMux I__9156 (
            .O(N__41089),
            .I(N__41081));
    LocalMux I__9155 (
            .O(N__41086),
            .I(N__41078));
    LocalMux I__9154 (
            .O(N__41081),
            .I(N__41075));
    Span4Mux_h I__9153 (
            .O(N__41078),
            .I(N__41069));
    Span4Mux_v I__9152 (
            .O(N__41075),
            .I(N__41066));
    InMux I__9151 (
            .O(N__41074),
            .I(N__41063));
    InMux I__9150 (
            .O(N__41073),
            .I(N__41058));
    InMux I__9149 (
            .O(N__41072),
            .I(N__41058));
    Span4Mux_v I__9148 (
            .O(N__41069),
            .I(N__41055));
    Span4Mux_h I__9147 (
            .O(N__41066),
            .I(N__41050));
    LocalMux I__9146 (
            .O(N__41063),
            .I(N__41050));
    LocalMux I__9145 (
            .O(N__41058),
            .I(N__41047));
    Odrv4 I__9144 (
            .O(N__41055),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__9143 (
            .O(N__41050),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__9142 (
            .O(N__41047),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__9141 (
            .O(N__41040),
            .I(N__41037));
    InMux I__9140 (
            .O(N__41037),
            .I(N__41034));
    LocalMux I__9139 (
            .O(N__41034),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__9138 (
            .O(N__41031),
            .I(N__41028));
    InMux I__9137 (
            .O(N__41028),
            .I(N__41025));
    LocalMux I__9136 (
            .O(N__41025),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__9135 (
            .O(N__41022),
            .I(N__41019));
    InMux I__9134 (
            .O(N__41019),
            .I(N__41016));
    LocalMux I__9133 (
            .O(N__41016),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ));
    InMux I__9132 (
            .O(N__41013),
            .I(N__41010));
    LocalMux I__9131 (
            .O(N__41010),
            .I(N__41007));
    Odrv4 I__9130 (
            .O(N__41007),
            .I(delay_hc_input_c));
    InMux I__9129 (
            .O(N__41004),
            .I(N__41001));
    LocalMux I__9128 (
            .O(N__41001),
            .I(N__40998));
    Span4Mux_h I__9127 (
            .O(N__40998),
            .I(N__40995));
    Span4Mux_v I__9126 (
            .O(N__40995),
            .I(N__40992));
    Odrv4 I__9125 (
            .O(N__40992),
            .I(delay_hc_d1));
    InMux I__9124 (
            .O(N__40989),
            .I(N__40985));
    InMux I__9123 (
            .O(N__40988),
            .I(N__40982));
    LocalMux I__9122 (
            .O(N__40985),
            .I(N__40979));
    LocalMux I__9121 (
            .O(N__40982),
            .I(N__40976));
    Span4Mux_v I__9120 (
            .O(N__40979),
            .I(N__40973));
    Span4Mux_v I__9119 (
            .O(N__40976),
            .I(N__40970));
    Span4Mux_v I__9118 (
            .O(N__40973),
            .I(N__40967));
    Span4Mux_h I__9117 (
            .O(N__40970),
            .I(N__40964));
    Odrv4 I__9116 (
            .O(N__40967),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__9115 (
            .O(N__40964),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__9114 (
            .O(N__40959),
            .I(N__40955));
    InMux I__9113 (
            .O(N__40958),
            .I(N__40951));
    LocalMux I__9112 (
            .O(N__40955),
            .I(N__40948));
    InMux I__9111 (
            .O(N__40954),
            .I(N__40945));
    LocalMux I__9110 (
            .O(N__40951),
            .I(N__40940));
    Span4Mux_h I__9109 (
            .O(N__40948),
            .I(N__40940));
    LocalMux I__9108 (
            .O(N__40945),
            .I(N__40937));
    Span4Mux_v I__9107 (
            .O(N__40940),
            .I(N__40934));
    Span4Mux_h I__9106 (
            .O(N__40937),
            .I(N__40931));
    Span4Mux_h I__9105 (
            .O(N__40934),
            .I(N__40928));
    Span4Mux_v I__9104 (
            .O(N__40931),
            .I(N__40925));
    Odrv4 I__9103 (
            .O(N__40928),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__9102 (
            .O(N__40925),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__9101 (
            .O(N__40920),
            .I(N__40917));
    LocalMux I__9100 (
            .O(N__40917),
            .I(N__40913));
    InMux I__9099 (
            .O(N__40916),
            .I(N__40908));
    Span4Mux_h I__9098 (
            .O(N__40913),
            .I(N__40905));
    InMux I__9097 (
            .O(N__40912),
            .I(N__40900));
    InMux I__9096 (
            .O(N__40911),
            .I(N__40900));
    LocalMux I__9095 (
            .O(N__40908),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    Odrv4 I__9094 (
            .O(N__40905),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    LocalMux I__9093 (
            .O(N__40900),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    InMux I__9092 (
            .O(N__40893),
            .I(N__40890));
    LocalMux I__9091 (
            .O(N__40890),
            .I(N__40887));
    Span4Mux_v I__9090 (
            .O(N__40887),
            .I(N__40882));
    InMux I__9089 (
            .O(N__40886),
            .I(N__40879));
    InMux I__9088 (
            .O(N__40885),
            .I(N__40874));
    Span4Mux_h I__9087 (
            .O(N__40882),
            .I(N__40871));
    LocalMux I__9086 (
            .O(N__40879),
            .I(N__40868));
    InMux I__9085 (
            .O(N__40878),
            .I(N__40865));
    InMux I__9084 (
            .O(N__40877),
            .I(N__40862));
    LocalMux I__9083 (
            .O(N__40874),
            .I(N__40859));
    Span4Mux_h I__9082 (
            .O(N__40871),
            .I(N__40854));
    Span4Mux_v I__9081 (
            .O(N__40868),
            .I(N__40854));
    LocalMux I__9080 (
            .O(N__40865),
            .I(N__40851));
    LocalMux I__9079 (
            .O(N__40862),
            .I(N__40844));
    Span4Mux_v I__9078 (
            .O(N__40859),
            .I(N__40844));
    Span4Mux_h I__9077 (
            .O(N__40854),
            .I(N__40844));
    Span4Mux_h I__9076 (
            .O(N__40851),
            .I(N__40841));
    Odrv4 I__9075 (
            .O(N__40844),
            .I(measured_delay_hc_2));
    Odrv4 I__9074 (
            .O(N__40841),
            .I(measured_delay_hc_2));
    InMux I__9073 (
            .O(N__40836),
            .I(N__40829));
    InMux I__9072 (
            .O(N__40835),
            .I(N__40824));
    InMux I__9071 (
            .O(N__40834),
            .I(N__40824));
    CascadeMux I__9070 (
            .O(N__40833),
            .I(N__40815));
    CascadeMux I__9069 (
            .O(N__40832),
            .I(N__40812));
    LocalMux I__9068 (
            .O(N__40829),
            .I(N__40803));
    LocalMux I__9067 (
            .O(N__40824),
            .I(N__40803));
    InMux I__9066 (
            .O(N__40823),
            .I(N__40795));
    InMux I__9065 (
            .O(N__40822),
            .I(N__40792));
    InMux I__9064 (
            .O(N__40821),
            .I(N__40787));
    InMux I__9063 (
            .O(N__40820),
            .I(N__40787));
    CascadeMux I__9062 (
            .O(N__40819),
            .I(N__40781));
    CascadeMux I__9061 (
            .O(N__40818),
            .I(N__40778));
    InMux I__9060 (
            .O(N__40815),
            .I(N__40770));
    InMux I__9059 (
            .O(N__40812),
            .I(N__40770));
    InMux I__9058 (
            .O(N__40811),
            .I(N__40763));
    InMux I__9057 (
            .O(N__40810),
            .I(N__40763));
    InMux I__9056 (
            .O(N__40809),
            .I(N__40763));
    InMux I__9055 (
            .O(N__40808),
            .I(N__40760));
    Span4Mux_h I__9054 (
            .O(N__40803),
            .I(N__40756));
    InMux I__9053 (
            .O(N__40802),
            .I(N__40753));
    InMux I__9052 (
            .O(N__40801),
            .I(N__40750));
    InMux I__9051 (
            .O(N__40800),
            .I(N__40745));
    InMux I__9050 (
            .O(N__40799),
            .I(N__40745));
    InMux I__9049 (
            .O(N__40798),
            .I(N__40737));
    LocalMux I__9048 (
            .O(N__40795),
            .I(N__40730));
    LocalMux I__9047 (
            .O(N__40792),
            .I(N__40730));
    LocalMux I__9046 (
            .O(N__40787),
            .I(N__40730));
    InMux I__9045 (
            .O(N__40786),
            .I(N__40723));
    InMux I__9044 (
            .O(N__40785),
            .I(N__40723));
    InMux I__9043 (
            .O(N__40784),
            .I(N__40723));
    InMux I__9042 (
            .O(N__40781),
            .I(N__40716));
    InMux I__9041 (
            .O(N__40778),
            .I(N__40716));
    InMux I__9040 (
            .O(N__40777),
            .I(N__40716));
    InMux I__9039 (
            .O(N__40776),
            .I(N__40711));
    InMux I__9038 (
            .O(N__40775),
            .I(N__40711));
    LocalMux I__9037 (
            .O(N__40770),
            .I(N__40706));
    LocalMux I__9036 (
            .O(N__40763),
            .I(N__40706));
    LocalMux I__9035 (
            .O(N__40760),
            .I(N__40703));
    InMux I__9034 (
            .O(N__40759),
            .I(N__40700));
    Sp12to4 I__9033 (
            .O(N__40756),
            .I(N__40691));
    LocalMux I__9032 (
            .O(N__40753),
            .I(N__40691));
    LocalMux I__9031 (
            .O(N__40750),
            .I(N__40691));
    LocalMux I__9030 (
            .O(N__40745),
            .I(N__40691));
    InMux I__9029 (
            .O(N__40744),
            .I(N__40684));
    InMux I__9028 (
            .O(N__40743),
            .I(N__40684));
    InMux I__9027 (
            .O(N__40742),
            .I(N__40684));
    InMux I__9026 (
            .O(N__40741),
            .I(N__40679));
    InMux I__9025 (
            .O(N__40740),
            .I(N__40679));
    LocalMux I__9024 (
            .O(N__40737),
            .I(N__40674));
    Span4Mux_v I__9023 (
            .O(N__40730),
            .I(N__40674));
    LocalMux I__9022 (
            .O(N__40723),
            .I(N__40665));
    LocalMux I__9021 (
            .O(N__40716),
            .I(N__40665));
    LocalMux I__9020 (
            .O(N__40711),
            .I(N__40665));
    Span4Mux_h I__9019 (
            .O(N__40706),
            .I(N__40665));
    Span4Mux_h I__9018 (
            .O(N__40703),
            .I(N__40662));
    LocalMux I__9017 (
            .O(N__40700),
            .I(N__40657));
    Span12Mux_v I__9016 (
            .O(N__40691),
            .I(N__40657));
    LocalMux I__9015 (
            .O(N__40684),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__9014 (
            .O(N__40679),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__9013 (
            .O(N__40674),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__9012 (
            .O(N__40665),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__9011 (
            .O(N__40662),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv12 I__9010 (
            .O(N__40657),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    InMux I__9009 (
            .O(N__40644),
            .I(N__40641));
    LocalMux I__9008 (
            .O(N__40641),
            .I(N__40636));
    InMux I__9007 (
            .O(N__40640),
            .I(N__40631));
    InMux I__9006 (
            .O(N__40639),
            .I(N__40631));
    Span4Mux_h I__9005 (
            .O(N__40636),
            .I(N__40614));
    LocalMux I__9004 (
            .O(N__40631),
            .I(N__40611));
    InMux I__9003 (
            .O(N__40630),
            .I(N__40604));
    InMux I__9002 (
            .O(N__40629),
            .I(N__40604));
    InMux I__9001 (
            .O(N__40628),
            .I(N__40604));
    InMux I__9000 (
            .O(N__40627),
            .I(N__40593));
    InMux I__8999 (
            .O(N__40626),
            .I(N__40593));
    InMux I__8998 (
            .O(N__40625),
            .I(N__40593));
    InMux I__8997 (
            .O(N__40624),
            .I(N__40593));
    InMux I__8996 (
            .O(N__40623),
            .I(N__40593));
    InMux I__8995 (
            .O(N__40622),
            .I(N__40590));
    InMux I__8994 (
            .O(N__40621),
            .I(N__40585));
    InMux I__8993 (
            .O(N__40620),
            .I(N__40585));
    InMux I__8992 (
            .O(N__40619),
            .I(N__40578));
    InMux I__8991 (
            .O(N__40618),
            .I(N__40578));
    InMux I__8990 (
            .O(N__40617),
            .I(N__40578));
    Odrv4 I__8989 (
            .O(N__40614),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv4 I__8988 (
            .O(N__40611),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__8987 (
            .O(N__40604),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__8986 (
            .O(N__40593),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__8985 (
            .O(N__40590),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__8984 (
            .O(N__40585),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__8983 (
            .O(N__40578),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    CascadeMux I__8982 (
            .O(N__40563),
            .I(N__40559));
    CascadeMux I__8981 (
            .O(N__40562),
            .I(N__40556));
    InMux I__8980 (
            .O(N__40559),
            .I(N__40551));
    InMux I__8979 (
            .O(N__40556),
            .I(N__40548));
    InMux I__8978 (
            .O(N__40555),
            .I(N__40545));
    InMux I__8977 (
            .O(N__40554),
            .I(N__40542));
    LocalMux I__8976 (
            .O(N__40551),
            .I(N__40537));
    LocalMux I__8975 (
            .O(N__40548),
            .I(N__40534));
    LocalMux I__8974 (
            .O(N__40545),
            .I(N__40531));
    LocalMux I__8973 (
            .O(N__40542),
            .I(N__40528));
    InMux I__8972 (
            .O(N__40541),
            .I(N__40525));
    CascadeMux I__8971 (
            .O(N__40540),
            .I(N__40522));
    Span4Mux_v I__8970 (
            .O(N__40537),
            .I(N__40519));
    Span4Mux_v I__8969 (
            .O(N__40534),
            .I(N__40514));
    Span4Mux_h I__8968 (
            .O(N__40531),
            .I(N__40514));
    Span4Mux_h I__8967 (
            .O(N__40528),
            .I(N__40511));
    LocalMux I__8966 (
            .O(N__40525),
            .I(N__40508));
    InMux I__8965 (
            .O(N__40522),
            .I(N__40505));
    Span4Mux_h I__8964 (
            .O(N__40519),
            .I(N__40500));
    Span4Mux_v I__8963 (
            .O(N__40514),
            .I(N__40500));
    Span4Mux_h I__8962 (
            .O(N__40511),
            .I(N__40497));
    Span12Mux_h I__8961 (
            .O(N__40508),
            .I(N__40494));
    LocalMux I__8960 (
            .O(N__40505),
            .I(measured_delay_hc_15));
    Odrv4 I__8959 (
            .O(N__40500),
            .I(measured_delay_hc_15));
    Odrv4 I__8958 (
            .O(N__40497),
            .I(measured_delay_hc_15));
    Odrv12 I__8957 (
            .O(N__40494),
            .I(measured_delay_hc_15));
    InMux I__8956 (
            .O(N__40485),
            .I(N__40481));
    InMux I__8955 (
            .O(N__40484),
            .I(N__40478));
    LocalMux I__8954 (
            .O(N__40481),
            .I(N__40475));
    LocalMux I__8953 (
            .O(N__40478),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv12 I__8952 (
            .O(N__40475),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__8951 (
            .O(N__40470),
            .I(N__40467));
    LocalMux I__8950 (
            .O(N__40467),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ));
    InMux I__8949 (
            .O(N__40464),
            .I(N__40460));
    InMux I__8948 (
            .O(N__40463),
            .I(N__40457));
    LocalMux I__8947 (
            .O(N__40460),
            .I(N__40454));
    LocalMux I__8946 (
            .O(N__40457),
            .I(N__40451));
    Odrv4 I__8945 (
            .O(N__40454),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__8944 (
            .O(N__40451),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__8943 (
            .O(N__40446),
            .I(N__40443));
    LocalMux I__8942 (
            .O(N__40443),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__8941 (
            .O(N__40440),
            .I(N__40437));
    InMux I__8940 (
            .O(N__40437),
            .I(N__40434));
    LocalMux I__8939 (
            .O(N__40434),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ));
    InMux I__8938 (
            .O(N__40431),
            .I(N__40428));
    LocalMux I__8937 (
            .O(N__40428),
            .I(N__40424));
    InMux I__8936 (
            .O(N__40427),
            .I(N__40421));
    Span4Mux_v I__8935 (
            .O(N__40424),
            .I(N__40416));
    LocalMux I__8934 (
            .O(N__40421),
            .I(N__40416));
    Odrv4 I__8933 (
            .O(N__40416),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__8932 (
            .O(N__40413),
            .I(N__40410));
    LocalMux I__8931 (
            .O(N__40410),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__8930 (
            .O(N__40407),
            .I(N__40404));
    InMux I__8929 (
            .O(N__40404),
            .I(N__40401));
    LocalMux I__8928 (
            .O(N__40401),
            .I(N__40398));
    Odrv4 I__8927 (
            .O(N__40398),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ));
    InMux I__8926 (
            .O(N__40395),
            .I(N__40392));
    LocalMux I__8925 (
            .O(N__40392),
            .I(N__40388));
    InMux I__8924 (
            .O(N__40391),
            .I(N__40385));
    Span4Mux_v I__8923 (
            .O(N__40388),
            .I(N__40380));
    LocalMux I__8922 (
            .O(N__40385),
            .I(N__40380));
    Odrv4 I__8921 (
            .O(N__40380),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__8920 (
            .O(N__40377),
            .I(N__40374));
    LocalMux I__8919 (
            .O(N__40374),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ));
    InMux I__8918 (
            .O(N__40371),
            .I(N__40368));
    LocalMux I__8917 (
            .O(N__40368),
            .I(N__40364));
    InMux I__8916 (
            .O(N__40367),
            .I(N__40361));
    Span4Mux_v I__8915 (
            .O(N__40364),
            .I(N__40358));
    LocalMux I__8914 (
            .O(N__40361),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__8913 (
            .O(N__40358),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__8912 (
            .O(N__40353),
            .I(N__40350));
    InMux I__8911 (
            .O(N__40350),
            .I(N__40347));
    LocalMux I__8910 (
            .O(N__40347),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ));
    InMux I__8909 (
            .O(N__40344),
            .I(N__40341));
    LocalMux I__8908 (
            .O(N__40341),
            .I(N__40337));
    InMux I__8907 (
            .O(N__40340),
            .I(N__40334));
    Span4Mux_v I__8906 (
            .O(N__40337),
            .I(N__40331));
    LocalMux I__8905 (
            .O(N__40334),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__8904 (
            .O(N__40331),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__8903 (
            .O(N__40326),
            .I(N__40323));
    LocalMux I__8902 (
            .O(N__40323),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ));
    InMux I__8901 (
            .O(N__40320),
            .I(N__40317));
    LocalMux I__8900 (
            .O(N__40317),
            .I(N__40313));
    InMux I__8899 (
            .O(N__40316),
            .I(N__40310));
    Span4Mux_v I__8898 (
            .O(N__40313),
            .I(N__40307));
    LocalMux I__8897 (
            .O(N__40310),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__8896 (
            .O(N__40307),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__8895 (
            .O(N__40302),
            .I(N__40299));
    LocalMux I__8894 (
            .O(N__40299),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ));
    InMux I__8893 (
            .O(N__40296),
            .I(N__40292));
    InMux I__8892 (
            .O(N__40295),
            .I(N__40289));
    LocalMux I__8891 (
            .O(N__40292),
            .I(N__40286));
    LocalMux I__8890 (
            .O(N__40289),
            .I(N__40283));
    Odrv4 I__8889 (
            .O(N__40286),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__8888 (
            .O(N__40283),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__8887 (
            .O(N__40278),
            .I(N__40275));
    LocalMux I__8886 (
            .O(N__40275),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__8885 (
            .O(N__40272),
            .I(N__40269));
    InMux I__8884 (
            .O(N__40269),
            .I(N__40266));
    LocalMux I__8883 (
            .O(N__40266),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ));
    InMux I__8882 (
            .O(N__40263),
            .I(N__40260));
    LocalMux I__8881 (
            .O(N__40260),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ));
    InMux I__8880 (
            .O(N__40257),
            .I(N__40254));
    LocalMux I__8879 (
            .O(N__40254),
            .I(N__40250));
    InMux I__8878 (
            .O(N__40253),
            .I(N__40247));
    Span4Mux_v I__8877 (
            .O(N__40250),
            .I(N__40242));
    LocalMux I__8876 (
            .O(N__40247),
            .I(N__40242));
    Odrv4 I__8875 (
            .O(N__40242),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__8874 (
            .O(N__40239),
            .I(N__40236));
    LocalMux I__8873 (
            .O(N__40236),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ));
    InMux I__8872 (
            .O(N__40233),
            .I(N__40229));
    InMux I__8871 (
            .O(N__40232),
            .I(N__40226));
    LocalMux I__8870 (
            .O(N__40229),
            .I(N__40223));
    LocalMux I__8869 (
            .O(N__40226),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__8868 (
            .O(N__40223),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__8867 (
            .O(N__40218),
            .I(N__40215));
    LocalMux I__8866 (
            .O(N__40215),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__8865 (
            .O(N__40212),
            .I(N__40209));
    InMux I__8864 (
            .O(N__40209),
            .I(N__40206));
    LocalMux I__8863 (
            .O(N__40206),
            .I(N__40203));
    Odrv4 I__8862 (
            .O(N__40203),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ));
    InMux I__8861 (
            .O(N__40200),
            .I(N__40197));
    LocalMux I__8860 (
            .O(N__40197),
            .I(N__40193));
    InMux I__8859 (
            .O(N__40196),
            .I(N__40190));
    Span4Mux_v I__8858 (
            .O(N__40193),
            .I(N__40187));
    LocalMux I__8857 (
            .O(N__40190),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__8856 (
            .O(N__40187),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__8855 (
            .O(N__40182),
            .I(N__40179));
    LocalMux I__8854 (
            .O(N__40179),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ));
    InMux I__8853 (
            .O(N__40176),
            .I(N__40172));
    InMux I__8852 (
            .O(N__40175),
            .I(N__40169));
    LocalMux I__8851 (
            .O(N__40172),
            .I(N__40166));
    LocalMux I__8850 (
            .O(N__40169),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv12 I__8849 (
            .O(N__40166),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__8848 (
            .O(N__40161),
            .I(N__40158));
    LocalMux I__8847 (
            .O(N__40158),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ));
    InMux I__8846 (
            .O(N__40155),
            .I(N__40151));
    InMux I__8845 (
            .O(N__40154),
            .I(N__40148));
    LocalMux I__8844 (
            .O(N__40151),
            .I(N__40145));
    LocalMux I__8843 (
            .O(N__40148),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv12 I__8842 (
            .O(N__40145),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__8841 (
            .O(N__40140),
            .I(N__40137));
    LocalMux I__8840 (
            .O(N__40137),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ));
    InMux I__8839 (
            .O(N__40134),
            .I(N__40130));
    InMux I__8838 (
            .O(N__40133),
            .I(N__40127));
    LocalMux I__8837 (
            .O(N__40130),
            .I(N__40124));
    LocalMux I__8836 (
            .O(N__40127),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv12 I__8835 (
            .O(N__40124),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__8834 (
            .O(N__40119),
            .I(N__40116));
    LocalMux I__8833 (
            .O(N__40116),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ));
    InMux I__8832 (
            .O(N__40113),
            .I(N__40109));
    InMux I__8831 (
            .O(N__40112),
            .I(N__40106));
    LocalMux I__8830 (
            .O(N__40109),
            .I(N__40103));
    LocalMux I__8829 (
            .O(N__40106),
            .I(N__40099));
    Span4Mux_h I__8828 (
            .O(N__40103),
            .I(N__40096));
    InMux I__8827 (
            .O(N__40102),
            .I(N__40093));
    Span4Mux_h I__8826 (
            .O(N__40099),
            .I(N__40090));
    Odrv4 I__8825 (
            .O(N__40096),
            .I(measured_delay_tr_2));
    LocalMux I__8824 (
            .O(N__40093),
            .I(measured_delay_tr_2));
    Odrv4 I__8823 (
            .O(N__40090),
            .I(measured_delay_tr_2));
    InMux I__8822 (
            .O(N__40083),
            .I(N__40080));
    LocalMux I__8821 (
            .O(N__40080),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ));
    InMux I__8820 (
            .O(N__40077),
            .I(N__40074));
    LocalMux I__8819 (
            .O(N__40074),
            .I(N__40070));
    CascadeMux I__8818 (
            .O(N__40073),
            .I(N__40067));
    Span4Mux_h I__8817 (
            .O(N__40070),
            .I(N__40064));
    InMux I__8816 (
            .O(N__40067),
            .I(N__40061));
    Odrv4 I__8815 (
            .O(N__40064),
            .I(measured_delay_tr_1));
    LocalMux I__8814 (
            .O(N__40061),
            .I(measured_delay_tr_1));
    CascadeMux I__8813 (
            .O(N__40056),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_ ));
    InMux I__8812 (
            .O(N__40053),
            .I(N__40050));
    LocalMux I__8811 (
            .O(N__40050),
            .I(N__40042));
    InMux I__8810 (
            .O(N__40049),
            .I(N__40037));
    InMux I__8809 (
            .O(N__40048),
            .I(N__40037));
    InMux I__8808 (
            .O(N__40047),
            .I(N__40030));
    InMux I__8807 (
            .O(N__40046),
            .I(N__40030));
    InMux I__8806 (
            .O(N__40045),
            .I(N__40030));
    Span4Mux_v I__8805 (
            .O(N__40042),
            .I(N__40025));
    LocalMux I__8804 (
            .O(N__40037),
            .I(N__40025));
    LocalMux I__8803 (
            .O(N__40030),
            .I(\phase_controller_inst1.stoper_tr.N_20_li ));
    Odrv4 I__8802 (
            .O(N__40025),
            .I(\phase_controller_inst1.stoper_tr.N_20_li ));
    CascadeMux I__8801 (
            .O(N__40020),
            .I(N__40016));
    CascadeMux I__8800 (
            .O(N__40019),
            .I(N__40011));
    InMux I__8799 (
            .O(N__40016),
            .I(N__40007));
    InMux I__8798 (
            .O(N__40015),
            .I(N__40002));
    InMux I__8797 (
            .O(N__40014),
            .I(N__40002));
    InMux I__8796 (
            .O(N__40011),
            .I(N__39999));
    InMux I__8795 (
            .O(N__40010),
            .I(N__39996));
    LocalMux I__8794 (
            .O(N__40007),
            .I(N__39991));
    LocalMux I__8793 (
            .O(N__40002),
            .I(N__39991));
    LocalMux I__8792 (
            .O(N__39999),
            .I(N__39984));
    LocalMux I__8791 (
            .O(N__39996),
            .I(N__39984));
    Span4Mux_v I__8790 (
            .O(N__39991),
            .I(N__39984));
    Odrv4 I__8789 (
            .O(N__39984),
            .I(measured_delay_tr_3));
    InMux I__8788 (
            .O(N__39981),
            .I(N__39978));
    LocalMux I__8787 (
            .O(N__39978),
            .I(N__39973));
    InMux I__8786 (
            .O(N__39977),
            .I(N__39969));
    InMux I__8785 (
            .O(N__39976),
            .I(N__39966));
    Span4Mux_v I__8784 (
            .O(N__39973),
            .I(N__39963));
    InMux I__8783 (
            .O(N__39972),
            .I(N__39960));
    LocalMux I__8782 (
            .O(N__39969),
            .I(N__39957));
    LocalMux I__8781 (
            .O(N__39966),
            .I(N__39952));
    Span4Mux_v I__8780 (
            .O(N__39963),
            .I(N__39952));
    LocalMux I__8779 (
            .O(N__39960),
            .I(N__39947));
    Span4Mux_h I__8778 (
            .O(N__39957),
            .I(N__39947));
    Odrv4 I__8777 (
            .O(N__39952),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__8776 (
            .O(N__39947),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__8775 (
            .O(N__39942),
            .I(N__39908));
    InMux I__8774 (
            .O(N__39941),
            .I(N__39908));
    InMux I__8773 (
            .O(N__39940),
            .I(N__39908));
    InMux I__8772 (
            .O(N__39939),
            .I(N__39908));
    InMux I__8771 (
            .O(N__39938),
            .I(N__39899));
    InMux I__8770 (
            .O(N__39937),
            .I(N__39899));
    InMux I__8769 (
            .O(N__39936),
            .I(N__39899));
    InMux I__8768 (
            .O(N__39935),
            .I(N__39899));
    InMux I__8767 (
            .O(N__39934),
            .I(N__39890));
    InMux I__8766 (
            .O(N__39933),
            .I(N__39890));
    InMux I__8765 (
            .O(N__39932),
            .I(N__39890));
    InMux I__8764 (
            .O(N__39931),
            .I(N__39890));
    InMux I__8763 (
            .O(N__39930),
            .I(N__39877));
    InMux I__8762 (
            .O(N__39929),
            .I(N__39877));
    InMux I__8761 (
            .O(N__39928),
            .I(N__39877));
    InMux I__8760 (
            .O(N__39927),
            .I(N__39877));
    InMux I__8759 (
            .O(N__39926),
            .I(N__39868));
    InMux I__8758 (
            .O(N__39925),
            .I(N__39868));
    InMux I__8757 (
            .O(N__39924),
            .I(N__39868));
    InMux I__8756 (
            .O(N__39923),
            .I(N__39868));
    InMux I__8755 (
            .O(N__39922),
            .I(N__39863));
    InMux I__8754 (
            .O(N__39921),
            .I(N__39863));
    InMux I__8753 (
            .O(N__39920),
            .I(N__39854));
    InMux I__8752 (
            .O(N__39919),
            .I(N__39854));
    InMux I__8751 (
            .O(N__39918),
            .I(N__39854));
    InMux I__8750 (
            .O(N__39917),
            .I(N__39854));
    LocalMux I__8749 (
            .O(N__39908),
            .I(N__39847));
    LocalMux I__8748 (
            .O(N__39899),
            .I(N__39847));
    LocalMux I__8747 (
            .O(N__39890),
            .I(N__39847));
    InMux I__8746 (
            .O(N__39889),
            .I(N__39838));
    InMux I__8745 (
            .O(N__39888),
            .I(N__39838));
    InMux I__8744 (
            .O(N__39887),
            .I(N__39838));
    InMux I__8743 (
            .O(N__39886),
            .I(N__39838));
    LocalMux I__8742 (
            .O(N__39877),
            .I(N__39835));
    LocalMux I__8741 (
            .O(N__39868),
            .I(N__39830));
    LocalMux I__8740 (
            .O(N__39863),
            .I(N__39830));
    LocalMux I__8739 (
            .O(N__39854),
            .I(N__39827));
    Span4Mux_v I__8738 (
            .O(N__39847),
            .I(N__39824));
    LocalMux I__8737 (
            .O(N__39838),
            .I(N__39815));
    Span4Mux_h I__8736 (
            .O(N__39835),
            .I(N__39815));
    Span4Mux_v I__8735 (
            .O(N__39830),
            .I(N__39815));
    Span4Mux_v I__8734 (
            .O(N__39827),
            .I(N__39815));
    Odrv4 I__8733 (
            .O(N__39824),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__8732 (
            .O(N__39815),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    CascadeMux I__8731 (
            .O(N__39810),
            .I(N__39807));
    InMux I__8730 (
            .O(N__39807),
            .I(N__39804));
    LocalMux I__8729 (
            .O(N__39804),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__8728 (
            .O(N__39801),
            .I(N__39798));
    InMux I__8727 (
            .O(N__39798),
            .I(N__39794));
    InMux I__8726 (
            .O(N__39797),
            .I(N__39790));
    LocalMux I__8725 (
            .O(N__39794),
            .I(N__39787));
    InMux I__8724 (
            .O(N__39793),
            .I(N__39784));
    LocalMux I__8723 (
            .O(N__39790),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__8722 (
            .O(N__39787),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__8721 (
            .O(N__39784),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__8720 (
            .O(N__39777),
            .I(N__39774));
    LocalMux I__8719 (
            .O(N__39774),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__8718 (
            .O(N__39771),
            .I(N__39768));
    InMux I__8717 (
            .O(N__39768),
            .I(N__39765));
    LocalMux I__8716 (
            .O(N__39765),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ));
    InMux I__8715 (
            .O(N__39762),
            .I(N__39758));
    InMux I__8714 (
            .O(N__39761),
            .I(N__39755));
    LocalMux I__8713 (
            .O(N__39758),
            .I(N__39752));
    LocalMux I__8712 (
            .O(N__39755),
            .I(N__39749));
    Odrv4 I__8711 (
            .O(N__39752),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__8710 (
            .O(N__39749),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__8709 (
            .O(N__39744),
            .I(N__39741));
    LocalMux I__8708 (
            .O(N__39741),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__8707 (
            .O(N__39738),
            .I(N__39735));
    InMux I__8706 (
            .O(N__39735),
            .I(N__39731));
    InMux I__8705 (
            .O(N__39734),
            .I(N__39728));
    LocalMux I__8704 (
            .O(N__39731),
            .I(N__39725));
    LocalMux I__8703 (
            .O(N__39728),
            .I(N__39722));
    Odrv4 I__8702 (
            .O(N__39725),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__8701 (
            .O(N__39722),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__8700 (
            .O(N__39717),
            .I(N__39714));
    InMux I__8699 (
            .O(N__39714),
            .I(N__39711));
    LocalMux I__8698 (
            .O(N__39711),
            .I(N__39708));
    Odrv4 I__8697 (
            .O(N__39708),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ));
    InMux I__8696 (
            .O(N__39705),
            .I(N__39702));
    LocalMux I__8695 (
            .O(N__39702),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ));
    InMux I__8694 (
            .O(N__39699),
            .I(N__39695));
    InMux I__8693 (
            .O(N__39698),
            .I(N__39692));
    LocalMux I__8692 (
            .O(N__39695),
            .I(N__39689));
    LocalMux I__8691 (
            .O(N__39692),
            .I(N__39686));
    Span4Mux_h I__8690 (
            .O(N__39689),
            .I(N__39683));
    Span4Mux_h I__8689 (
            .O(N__39686),
            .I(N__39680));
    Odrv4 I__8688 (
            .O(N__39683),
            .I(\delay_measurement_inst.N_284_1 ));
    Odrv4 I__8687 (
            .O(N__39680),
            .I(\delay_measurement_inst.N_284_1 ));
    InMux I__8686 (
            .O(N__39675),
            .I(N__39672));
    LocalMux I__8685 (
            .O(N__39672),
            .I(N__39666));
    InMux I__8684 (
            .O(N__39671),
            .I(N__39662));
    InMux I__8683 (
            .O(N__39670),
            .I(N__39657));
    InMux I__8682 (
            .O(N__39669),
            .I(N__39657));
    Span4Mux_h I__8681 (
            .O(N__39666),
            .I(N__39654));
    InMux I__8680 (
            .O(N__39665),
            .I(N__39650));
    LocalMux I__8679 (
            .O(N__39662),
            .I(N__39647));
    LocalMux I__8678 (
            .O(N__39657),
            .I(N__39644));
    Span4Mux_v I__8677 (
            .O(N__39654),
            .I(N__39640));
    InMux I__8676 (
            .O(N__39653),
            .I(N__39637));
    LocalMux I__8675 (
            .O(N__39650),
            .I(N__39630));
    Span4Mux_v I__8674 (
            .O(N__39647),
            .I(N__39630));
    Span4Mux_h I__8673 (
            .O(N__39644),
            .I(N__39630));
    InMux I__8672 (
            .O(N__39643),
            .I(N__39627));
    Odrv4 I__8671 (
            .O(N__39640),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    LocalMux I__8670 (
            .O(N__39637),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    Odrv4 I__8669 (
            .O(N__39630),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    LocalMux I__8668 (
            .O(N__39627),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    InMux I__8667 (
            .O(N__39618),
            .I(N__39615));
    LocalMux I__8666 (
            .O(N__39615),
            .I(N__39611));
    InMux I__8665 (
            .O(N__39614),
            .I(N__39608));
    Span4Mux_v I__8664 (
            .O(N__39611),
            .I(N__39603));
    LocalMux I__8663 (
            .O(N__39608),
            .I(N__39603));
    Span4Mux_h I__8662 (
            .O(N__39603),
            .I(N__39599));
    InMux I__8661 (
            .O(N__39602),
            .I(N__39596));
    Odrv4 I__8660 (
            .O(N__39599),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i ));
    LocalMux I__8659 (
            .O(N__39596),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i ));
    InMux I__8658 (
            .O(N__39591),
            .I(N__39588));
    LocalMux I__8657 (
            .O(N__39588),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ));
    InMux I__8656 (
            .O(N__39585),
            .I(N__39582));
    LocalMux I__8655 (
            .O(N__39582),
            .I(N__39579));
    Span4Mux_v I__8654 (
            .O(N__39579),
            .I(N__39576));
    Span4Mux_h I__8653 (
            .O(N__39576),
            .I(N__39571));
    InMux I__8652 (
            .O(N__39575),
            .I(N__39568));
    InMux I__8651 (
            .O(N__39574),
            .I(N__39565));
    Odrv4 I__8650 (
            .O(N__39571),
            .I(measured_delay_tr_8));
    LocalMux I__8649 (
            .O(N__39568),
            .I(measured_delay_tr_8));
    LocalMux I__8648 (
            .O(N__39565),
            .I(measured_delay_tr_8));
    InMux I__8647 (
            .O(N__39558),
            .I(N__39555));
    LocalMux I__8646 (
            .O(N__39555),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ));
    InMux I__8645 (
            .O(N__39552),
            .I(N__39549));
    LocalMux I__8644 (
            .O(N__39549),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ));
    InMux I__8643 (
            .O(N__39546),
            .I(N__39543));
    LocalMux I__8642 (
            .O(N__39543),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ));
    InMux I__8641 (
            .O(N__39540),
            .I(N__39537));
    LocalMux I__8640 (
            .O(N__39537),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    InMux I__8639 (
            .O(N__39534),
            .I(N__39531));
    LocalMux I__8638 (
            .O(N__39531),
            .I(N__39525));
    InMux I__8637 (
            .O(N__39530),
            .I(N__39520));
    InMux I__8636 (
            .O(N__39529),
            .I(N__39520));
    InMux I__8635 (
            .O(N__39528),
            .I(N__39517));
    Span4Mux_h I__8634 (
            .O(N__39525),
            .I(N__39514));
    LocalMux I__8633 (
            .O(N__39520),
            .I(N__39511));
    LocalMux I__8632 (
            .O(N__39517),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    Odrv4 I__8631 (
            .O(N__39514),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    Odrv12 I__8630 (
            .O(N__39511),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    InMux I__8629 (
            .O(N__39504),
            .I(N__39501));
    LocalMux I__8628 (
            .O(N__39501),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ));
    InMux I__8627 (
            .O(N__39498),
            .I(N__39495));
    LocalMux I__8626 (
            .O(N__39495),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ));
    InMux I__8625 (
            .O(N__39492),
            .I(N__39489));
    LocalMux I__8624 (
            .O(N__39489),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ));
    InMux I__8623 (
            .O(N__39486),
            .I(N__39483));
    LocalMux I__8622 (
            .O(N__39483),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ));
    CascadeMux I__8621 (
            .O(N__39480),
            .I(N__39477));
    InMux I__8620 (
            .O(N__39477),
            .I(N__39474));
    LocalMux I__8619 (
            .O(N__39474),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ));
    InMux I__8618 (
            .O(N__39471),
            .I(N__39468));
    LocalMux I__8617 (
            .O(N__39468),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__8616 (
            .O(N__39465),
            .I(N__39462));
    InMux I__8615 (
            .O(N__39462),
            .I(N__39459));
    LocalMux I__8614 (
            .O(N__39459),
            .I(N__39456));
    Odrv4 I__8613 (
            .O(N__39456),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ));
    InMux I__8612 (
            .O(N__39453),
            .I(N__39450));
    LocalMux I__8611 (
            .O(N__39450),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__8610 (
            .O(N__39447),
            .I(N__39444));
    InMux I__8609 (
            .O(N__39444),
            .I(N__39441));
    LocalMux I__8608 (
            .O(N__39441),
            .I(N__39438));
    Span4Mux_h I__8607 (
            .O(N__39438),
            .I(N__39435));
    Odrv4 I__8606 (
            .O(N__39435),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ));
    InMux I__8605 (
            .O(N__39432),
            .I(N__39429));
    LocalMux I__8604 (
            .O(N__39429),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ));
    CascadeMux I__8603 (
            .O(N__39426),
            .I(N__39423));
    InMux I__8602 (
            .O(N__39423),
            .I(N__39420));
    LocalMux I__8601 (
            .O(N__39420),
            .I(N__39417));
    Span4Mux_h I__8600 (
            .O(N__39417),
            .I(N__39414));
    Odrv4 I__8599 (
            .O(N__39414),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ));
    InMux I__8598 (
            .O(N__39411),
            .I(N__39408));
    LocalMux I__8597 (
            .O(N__39408),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ));
    CascadeMux I__8596 (
            .O(N__39405),
            .I(N__39402));
    InMux I__8595 (
            .O(N__39402),
            .I(N__39399));
    LocalMux I__8594 (
            .O(N__39399),
            .I(N__39396));
    Span4Mux_h I__8593 (
            .O(N__39396),
            .I(N__39393));
    Odrv4 I__8592 (
            .O(N__39393),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ));
    InMux I__8591 (
            .O(N__39390),
            .I(N__39387));
    LocalMux I__8590 (
            .O(N__39387),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ));
    InMux I__8589 (
            .O(N__39384),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__8588 (
            .O(N__39381),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ));
    InMux I__8587 (
            .O(N__39378),
            .I(N__39375));
    LocalMux I__8586 (
            .O(N__39375),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__8585 (
            .O(N__39372),
            .I(N__39369));
    InMux I__8584 (
            .O(N__39369),
            .I(N__39366));
    LocalMux I__8583 (
            .O(N__39366),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ));
    InMux I__8582 (
            .O(N__39363),
            .I(N__39360));
    LocalMux I__8581 (
            .O(N__39360),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__8580 (
            .O(N__39357),
            .I(N__39354));
    InMux I__8579 (
            .O(N__39354),
            .I(N__39351));
    LocalMux I__8578 (
            .O(N__39351),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ));
    InMux I__8577 (
            .O(N__39348),
            .I(N__39345));
    LocalMux I__8576 (
            .O(N__39345),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__8575 (
            .O(N__39342),
            .I(N__39339));
    InMux I__8574 (
            .O(N__39339),
            .I(N__39336));
    LocalMux I__8573 (
            .O(N__39336),
            .I(N__39333));
    Odrv12 I__8572 (
            .O(N__39333),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ));
    InMux I__8571 (
            .O(N__39330),
            .I(N__39327));
    LocalMux I__8570 (
            .O(N__39327),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__8569 (
            .O(N__39324),
            .I(N__39321));
    InMux I__8568 (
            .O(N__39321),
            .I(N__39318));
    LocalMux I__8567 (
            .O(N__39318),
            .I(N__39315));
    Odrv4 I__8566 (
            .O(N__39315),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ));
    InMux I__8565 (
            .O(N__39312),
            .I(N__39309));
    LocalMux I__8564 (
            .O(N__39309),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__8563 (
            .O(N__39306),
            .I(N__39303));
    InMux I__8562 (
            .O(N__39303),
            .I(N__39300));
    LocalMux I__8561 (
            .O(N__39300),
            .I(N__39297));
    Span4Mux_h I__8560 (
            .O(N__39297),
            .I(N__39294));
    Span4Mux_h I__8559 (
            .O(N__39294),
            .I(N__39291));
    Odrv4 I__8558 (
            .O(N__39291),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ));
    InMux I__8557 (
            .O(N__39288),
            .I(N__39285));
    LocalMux I__8556 (
            .O(N__39285),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__8555 (
            .O(N__39282),
            .I(N__39279));
    InMux I__8554 (
            .O(N__39279),
            .I(N__39276));
    LocalMux I__8553 (
            .O(N__39276),
            .I(N__39273));
    Span4Mux_h I__8552 (
            .O(N__39273),
            .I(N__39270));
    Odrv4 I__8551 (
            .O(N__39270),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ));
    InMux I__8550 (
            .O(N__39267),
            .I(N__39264));
    LocalMux I__8549 (
            .O(N__39264),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ));
    InMux I__8548 (
            .O(N__39261),
            .I(N__39258));
    LocalMux I__8547 (
            .O(N__39258),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__8546 (
            .O(N__39255),
            .I(N__39252));
    InMux I__8545 (
            .O(N__39252),
            .I(N__39249));
    LocalMux I__8544 (
            .O(N__39249),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__8543 (
            .O(N__39246),
            .I(N__39243));
    InMux I__8542 (
            .O(N__39243),
            .I(N__39240));
    LocalMux I__8541 (
            .O(N__39240),
            .I(N__39237));
    Odrv4 I__8540 (
            .O(N__39237),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ));
    InMux I__8539 (
            .O(N__39234),
            .I(N__39231));
    LocalMux I__8538 (
            .O(N__39231),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ));
    InMux I__8537 (
            .O(N__39228),
            .I(N__39225));
    LocalMux I__8536 (
            .O(N__39225),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ));
    InMux I__8535 (
            .O(N__39222),
            .I(N__39219));
    LocalMux I__8534 (
            .O(N__39219),
            .I(N__39216));
    Odrv12 I__8533 (
            .O(N__39216),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_6 ));
    CascadeMux I__8532 (
            .O(N__39213),
            .I(N__39210));
    InMux I__8531 (
            .O(N__39210),
            .I(N__39207));
    LocalMux I__8530 (
            .O(N__39207),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__8529 (
            .O(N__39204),
            .I(N__39201));
    InMux I__8528 (
            .O(N__39201),
            .I(N__39198));
    LocalMux I__8527 (
            .O(N__39198),
            .I(N__39195));
    Odrv4 I__8526 (
            .O(N__39195),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ));
    InMux I__8525 (
            .O(N__39192),
            .I(N__39189));
    LocalMux I__8524 (
            .O(N__39189),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__8523 (
            .O(N__39186),
            .I(N__39183));
    InMux I__8522 (
            .O(N__39183),
            .I(N__39180));
    LocalMux I__8521 (
            .O(N__39180),
            .I(N__39177));
    Odrv4 I__8520 (
            .O(N__39177),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ));
    InMux I__8519 (
            .O(N__39174),
            .I(N__39171));
    LocalMux I__8518 (
            .O(N__39171),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__8517 (
            .O(N__39168),
            .I(N__39165));
    InMux I__8516 (
            .O(N__39165),
            .I(N__39162));
    LocalMux I__8515 (
            .O(N__39162),
            .I(N__39159));
    Odrv4 I__8514 (
            .O(N__39159),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ));
    InMux I__8513 (
            .O(N__39156),
            .I(N__39153));
    LocalMux I__8512 (
            .O(N__39153),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__8511 (
            .O(N__39150),
            .I(N__39147));
    InMux I__8510 (
            .O(N__39147),
            .I(N__39144));
    LocalMux I__8509 (
            .O(N__39144),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ));
    InMux I__8508 (
            .O(N__39141),
            .I(N__39138));
    LocalMux I__8507 (
            .O(N__39138),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__8506 (
            .O(N__39135),
            .I(N__39132));
    InMux I__8505 (
            .O(N__39132),
            .I(N__39129));
    LocalMux I__8504 (
            .O(N__39129),
            .I(N__39126));
    Odrv4 I__8503 (
            .O(N__39126),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ));
    InMux I__8502 (
            .O(N__39123),
            .I(N__39120));
    LocalMux I__8501 (
            .O(N__39120),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__8500 (
            .O(N__39117),
            .I(N__39114));
    InMux I__8499 (
            .O(N__39114),
            .I(N__39111));
    LocalMux I__8498 (
            .O(N__39111),
            .I(N__39108));
    Odrv4 I__8497 (
            .O(N__39108),
            .I(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ));
    InMux I__8496 (
            .O(N__39105),
            .I(N__39102));
    LocalMux I__8495 (
            .O(N__39102),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__8494 (
            .O(N__39099),
            .I(N__39096));
    InMux I__8493 (
            .O(N__39096),
            .I(N__39093));
    LocalMux I__8492 (
            .O(N__39093),
            .I(N__39090));
    Odrv4 I__8491 (
            .O(N__39090),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ));
    CascadeMux I__8490 (
            .O(N__39087),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_ ));
    InMux I__8489 (
            .O(N__39084),
            .I(N__39081));
    LocalMux I__8488 (
            .O(N__39081),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0 ));
    InMux I__8487 (
            .O(N__39078),
            .I(N__39074));
    InMux I__8486 (
            .O(N__39077),
            .I(N__39071));
    LocalMux I__8485 (
            .O(N__39074),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    LocalMux I__8484 (
            .O(N__39071),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    InMux I__8483 (
            .O(N__39066),
            .I(N__39063));
    LocalMux I__8482 (
            .O(N__39063),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_0 ));
    InMux I__8481 (
            .O(N__39060),
            .I(N__39057));
    LocalMux I__8480 (
            .O(N__39057),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4 ));
    CascadeMux I__8479 (
            .O(N__39054),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_ ));
    InMux I__8478 (
            .O(N__39051),
            .I(N__39048));
    LocalMux I__8477 (
            .O(N__39048),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ));
    CascadeMux I__8476 (
            .O(N__39045),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_cascade_ ));
    InMux I__8475 (
            .O(N__39042),
            .I(N__39034));
    InMux I__8474 (
            .O(N__39041),
            .I(N__39031));
    InMux I__8473 (
            .O(N__39040),
            .I(N__39022));
    InMux I__8472 (
            .O(N__39039),
            .I(N__39022));
    InMux I__8471 (
            .O(N__39038),
            .I(N__39019));
    InMux I__8470 (
            .O(N__39037),
            .I(N__39016));
    LocalMux I__8469 (
            .O(N__39034),
            .I(N__39010));
    LocalMux I__8468 (
            .O(N__39031),
            .I(N__39010));
    InMux I__8467 (
            .O(N__39030),
            .I(N__39007));
    InMux I__8466 (
            .O(N__39029),
            .I(N__38998));
    InMux I__8465 (
            .O(N__39028),
            .I(N__38998));
    InMux I__8464 (
            .O(N__39027),
            .I(N__38998));
    LocalMux I__8463 (
            .O(N__39022),
            .I(N__38995));
    LocalMux I__8462 (
            .O(N__39019),
            .I(N__38990));
    LocalMux I__8461 (
            .O(N__39016),
            .I(N__38990));
    InMux I__8460 (
            .O(N__39015),
            .I(N__38987));
    Span4Mux_h I__8459 (
            .O(N__39010),
            .I(N__38982));
    LocalMux I__8458 (
            .O(N__39007),
            .I(N__38982));
    InMux I__8457 (
            .O(N__39006),
            .I(N__38979));
    InMux I__8456 (
            .O(N__39005),
            .I(N__38976));
    LocalMux I__8455 (
            .O(N__38998),
            .I(N__38973));
    Span4Mux_v I__8454 (
            .O(N__38995),
            .I(N__38966));
    Span4Mux_v I__8453 (
            .O(N__38990),
            .I(N__38966));
    LocalMux I__8452 (
            .O(N__38987),
            .I(N__38966));
    Span4Mux_h I__8451 (
            .O(N__38982),
            .I(N__38961));
    LocalMux I__8450 (
            .O(N__38979),
            .I(N__38961));
    LocalMux I__8449 (
            .O(N__38976),
            .I(N__38958));
    Span4Mux_v I__8448 (
            .O(N__38973),
            .I(N__38955));
    Span4Mux_h I__8447 (
            .O(N__38966),
            .I(N__38948));
    Span4Mux_v I__8446 (
            .O(N__38961),
            .I(N__38948));
    Span4Mux_v I__8445 (
            .O(N__38958),
            .I(N__38948));
    Odrv4 I__8444 (
            .O(N__38955),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    Odrv4 I__8443 (
            .O(N__38948),
            .I(\delay_measurement_inst.delay_hc_reg3lt31_0 ));
    InMux I__8442 (
            .O(N__38943),
            .I(N__38940));
    LocalMux I__8441 (
            .O(N__38940),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4 ));
    CascadeMux I__8440 (
            .O(N__38937),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_5_cascade_ ));
    CascadeMux I__8439 (
            .O(N__38934),
            .I(N__38931));
    InMux I__8438 (
            .O(N__38931),
            .I(N__38928));
    LocalMux I__8437 (
            .O(N__38928),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0 ));
    InMux I__8436 (
            .O(N__38925),
            .I(N__38922));
    LocalMux I__8435 (
            .O(N__38922),
            .I(N__38919));
    Odrv4 I__8434 (
            .O(N__38919),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19 ));
    CascadeMux I__8433 (
            .O(N__38916),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_ ));
    InMux I__8432 (
            .O(N__38913),
            .I(N__38910));
    LocalMux I__8431 (
            .O(N__38910),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ));
    InMux I__8430 (
            .O(N__38907),
            .I(N__38904));
    LocalMux I__8429 (
            .O(N__38904),
            .I(N__38901));
    Odrv4 I__8428 (
            .O(N__38901),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0 ));
    InMux I__8427 (
            .O(N__38898),
            .I(N__38895));
    LocalMux I__8426 (
            .O(N__38895),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7 ));
    InMux I__8425 (
            .O(N__38892),
            .I(N__38889));
    LocalMux I__8424 (
            .O(N__38889),
            .I(N__38886));
    Odrv4 I__8423 (
            .O(N__38886),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3 ));
    InMux I__8422 (
            .O(N__38883),
            .I(N__38880));
    LocalMux I__8421 (
            .O(N__38880),
            .I(N__38877));
    Odrv4 I__8420 (
            .O(N__38877),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1 ));
    CascadeMux I__8419 (
            .O(N__38874),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz_cascade_ ));
    CascadeMux I__8418 (
            .O(N__38871),
            .I(N__38866));
    InMux I__8417 (
            .O(N__38870),
            .I(N__38863));
    InMux I__8416 (
            .O(N__38869),
            .I(N__38860));
    InMux I__8415 (
            .O(N__38866),
            .I(N__38857));
    LocalMux I__8414 (
            .O(N__38863),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__8413 (
            .O(N__38860),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__8412 (
            .O(N__38857),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__8411 (
            .O(N__38850),
            .I(bfn_15_22_0_));
    CascadeMux I__8410 (
            .O(N__38847),
            .I(N__38842));
    InMux I__8409 (
            .O(N__38846),
            .I(N__38839));
    InMux I__8408 (
            .O(N__38845),
            .I(N__38836));
    InMux I__8407 (
            .O(N__38842),
            .I(N__38833));
    LocalMux I__8406 (
            .O(N__38839),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__8405 (
            .O(N__38836),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__8404 (
            .O(N__38833),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__8403 (
            .O(N__38826),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    CascadeMux I__8402 (
            .O(N__38823),
            .I(N__38818));
    InMux I__8401 (
            .O(N__38822),
            .I(N__38815));
    InMux I__8400 (
            .O(N__38821),
            .I(N__38812));
    InMux I__8399 (
            .O(N__38818),
            .I(N__38809));
    LocalMux I__8398 (
            .O(N__38815),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__8397 (
            .O(N__38812),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__8396 (
            .O(N__38809),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__8395 (
            .O(N__38802),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    CascadeMux I__8394 (
            .O(N__38799),
            .I(N__38794));
    InMux I__8393 (
            .O(N__38798),
            .I(N__38791));
    InMux I__8392 (
            .O(N__38797),
            .I(N__38788));
    InMux I__8391 (
            .O(N__38794),
            .I(N__38785));
    LocalMux I__8390 (
            .O(N__38791),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__8389 (
            .O(N__38788),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__8388 (
            .O(N__38785),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__8387 (
            .O(N__38778),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    CascadeMux I__8386 (
            .O(N__38775),
            .I(N__38771));
    InMux I__8385 (
            .O(N__38774),
            .I(N__38768));
    InMux I__8384 (
            .O(N__38771),
            .I(N__38765));
    LocalMux I__8383 (
            .O(N__38768),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__8382 (
            .O(N__38765),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__8381 (
            .O(N__38760),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__8380 (
            .O(N__38757),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CascadeMux I__8379 (
            .O(N__38754),
            .I(N__38750));
    InMux I__8378 (
            .O(N__38753),
            .I(N__38747));
    InMux I__8377 (
            .O(N__38750),
            .I(N__38744));
    LocalMux I__8376 (
            .O(N__38747),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__8375 (
            .O(N__38744),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__8374 (
            .O(N__38739),
            .I(N__38736));
    LocalMux I__8373 (
            .O(N__38736),
            .I(N__38733));
    Span4Mux_v I__8372 (
            .O(N__38733),
            .I(N__38728));
    CEMux I__8371 (
            .O(N__38732),
            .I(N__38725));
    CEMux I__8370 (
            .O(N__38731),
            .I(N__38721));
    Span4Mux_h I__8369 (
            .O(N__38728),
            .I(N__38716));
    LocalMux I__8368 (
            .O(N__38725),
            .I(N__38716));
    CEMux I__8367 (
            .O(N__38724),
            .I(N__38713));
    LocalMux I__8366 (
            .O(N__38721),
            .I(N__38710));
    Span4Mux_v I__8365 (
            .O(N__38716),
            .I(N__38707));
    LocalMux I__8364 (
            .O(N__38713),
            .I(N__38702));
    Span4Mux_v I__8363 (
            .O(N__38710),
            .I(N__38702));
    Odrv4 I__8362 (
            .O(N__38707),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    Odrv4 I__8361 (
            .O(N__38702),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    CascadeMux I__8360 (
            .O(N__38697),
            .I(N__38692));
    InMux I__8359 (
            .O(N__38696),
            .I(N__38689));
    InMux I__8358 (
            .O(N__38695),
            .I(N__38686));
    InMux I__8357 (
            .O(N__38692),
            .I(N__38683));
    LocalMux I__8356 (
            .O(N__38689),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__8355 (
            .O(N__38686),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__8354 (
            .O(N__38683),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__8353 (
            .O(N__38676),
            .I(bfn_15_21_0_));
    CascadeMux I__8352 (
            .O(N__38673),
            .I(N__38668));
    InMux I__8351 (
            .O(N__38672),
            .I(N__38665));
    InMux I__8350 (
            .O(N__38671),
            .I(N__38662));
    InMux I__8349 (
            .O(N__38668),
            .I(N__38659));
    LocalMux I__8348 (
            .O(N__38665),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__8347 (
            .O(N__38662),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__8346 (
            .O(N__38659),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__8345 (
            .O(N__38652),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    CascadeMux I__8344 (
            .O(N__38649),
            .I(N__38644));
    InMux I__8343 (
            .O(N__38648),
            .I(N__38641));
    InMux I__8342 (
            .O(N__38647),
            .I(N__38638));
    InMux I__8341 (
            .O(N__38644),
            .I(N__38635));
    LocalMux I__8340 (
            .O(N__38641),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__8339 (
            .O(N__38638),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__8338 (
            .O(N__38635),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__8337 (
            .O(N__38628),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    CascadeMux I__8336 (
            .O(N__38625),
            .I(N__38620));
    InMux I__8335 (
            .O(N__38624),
            .I(N__38617));
    InMux I__8334 (
            .O(N__38623),
            .I(N__38614));
    InMux I__8333 (
            .O(N__38620),
            .I(N__38611));
    LocalMux I__8332 (
            .O(N__38617),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__8331 (
            .O(N__38614),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__8330 (
            .O(N__38611),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__8329 (
            .O(N__38604),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    CascadeMux I__8328 (
            .O(N__38601),
            .I(N__38596));
    InMux I__8327 (
            .O(N__38600),
            .I(N__38593));
    InMux I__8326 (
            .O(N__38599),
            .I(N__38590));
    InMux I__8325 (
            .O(N__38596),
            .I(N__38587));
    LocalMux I__8324 (
            .O(N__38593),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__8323 (
            .O(N__38590),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__8322 (
            .O(N__38587),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__8321 (
            .O(N__38580),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    CascadeMux I__8320 (
            .O(N__38577),
            .I(N__38572));
    InMux I__8319 (
            .O(N__38576),
            .I(N__38569));
    InMux I__8318 (
            .O(N__38575),
            .I(N__38566));
    InMux I__8317 (
            .O(N__38572),
            .I(N__38563));
    LocalMux I__8316 (
            .O(N__38569),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__8315 (
            .O(N__38566),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__8314 (
            .O(N__38563),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__8313 (
            .O(N__38556),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    CascadeMux I__8312 (
            .O(N__38553),
            .I(N__38548));
    InMux I__8311 (
            .O(N__38552),
            .I(N__38545));
    InMux I__8310 (
            .O(N__38551),
            .I(N__38542));
    InMux I__8309 (
            .O(N__38548),
            .I(N__38539));
    LocalMux I__8308 (
            .O(N__38545),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__8307 (
            .O(N__38542),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__8306 (
            .O(N__38539),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__8305 (
            .O(N__38532),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    CascadeMux I__8304 (
            .O(N__38529),
            .I(N__38524));
    InMux I__8303 (
            .O(N__38528),
            .I(N__38521));
    InMux I__8302 (
            .O(N__38527),
            .I(N__38518));
    InMux I__8301 (
            .O(N__38524),
            .I(N__38515));
    LocalMux I__8300 (
            .O(N__38521),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__8299 (
            .O(N__38518),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__8298 (
            .O(N__38515),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__8297 (
            .O(N__38508),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    CascadeMux I__8296 (
            .O(N__38505),
            .I(N__38500));
    InMux I__8295 (
            .O(N__38504),
            .I(N__38497));
    InMux I__8294 (
            .O(N__38503),
            .I(N__38494));
    InMux I__8293 (
            .O(N__38500),
            .I(N__38491));
    LocalMux I__8292 (
            .O(N__38497),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__8291 (
            .O(N__38494),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__8290 (
            .O(N__38491),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__8289 (
            .O(N__38484),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    CascadeMux I__8288 (
            .O(N__38481),
            .I(N__38476));
    InMux I__8287 (
            .O(N__38480),
            .I(N__38473));
    InMux I__8286 (
            .O(N__38479),
            .I(N__38470));
    InMux I__8285 (
            .O(N__38476),
            .I(N__38467));
    LocalMux I__8284 (
            .O(N__38473),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__8283 (
            .O(N__38470),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__8282 (
            .O(N__38467),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__8281 (
            .O(N__38460),
            .I(bfn_15_20_0_));
    CascadeMux I__8280 (
            .O(N__38457),
            .I(N__38452));
    InMux I__8279 (
            .O(N__38456),
            .I(N__38449));
    InMux I__8278 (
            .O(N__38455),
            .I(N__38446));
    InMux I__8277 (
            .O(N__38452),
            .I(N__38443));
    LocalMux I__8276 (
            .O(N__38449),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__8275 (
            .O(N__38446),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__8274 (
            .O(N__38443),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__8273 (
            .O(N__38436),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__8272 (
            .O(N__38433),
            .I(N__38428));
    InMux I__8271 (
            .O(N__38432),
            .I(N__38425));
    InMux I__8270 (
            .O(N__38431),
            .I(N__38422));
    InMux I__8269 (
            .O(N__38428),
            .I(N__38419));
    LocalMux I__8268 (
            .O(N__38425),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__8267 (
            .O(N__38422),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__8266 (
            .O(N__38419),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__8265 (
            .O(N__38412),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    CascadeMux I__8264 (
            .O(N__38409),
            .I(N__38404));
    InMux I__8263 (
            .O(N__38408),
            .I(N__38401));
    InMux I__8262 (
            .O(N__38407),
            .I(N__38398));
    InMux I__8261 (
            .O(N__38404),
            .I(N__38395));
    LocalMux I__8260 (
            .O(N__38401),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__8259 (
            .O(N__38398),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__8258 (
            .O(N__38395),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__8257 (
            .O(N__38388),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    CascadeMux I__8256 (
            .O(N__38385),
            .I(N__38380));
    InMux I__8255 (
            .O(N__38384),
            .I(N__38377));
    InMux I__8254 (
            .O(N__38383),
            .I(N__38374));
    InMux I__8253 (
            .O(N__38380),
            .I(N__38371));
    LocalMux I__8252 (
            .O(N__38377),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__8251 (
            .O(N__38374),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__8250 (
            .O(N__38371),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__8249 (
            .O(N__38364),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    CascadeMux I__8248 (
            .O(N__38361),
            .I(N__38356));
    InMux I__8247 (
            .O(N__38360),
            .I(N__38353));
    InMux I__8246 (
            .O(N__38359),
            .I(N__38350));
    InMux I__8245 (
            .O(N__38356),
            .I(N__38347));
    LocalMux I__8244 (
            .O(N__38353),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__8243 (
            .O(N__38350),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__8242 (
            .O(N__38347),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__8241 (
            .O(N__38340),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    CascadeMux I__8240 (
            .O(N__38337),
            .I(N__38332));
    InMux I__8239 (
            .O(N__38336),
            .I(N__38329));
    InMux I__8238 (
            .O(N__38335),
            .I(N__38326));
    InMux I__8237 (
            .O(N__38332),
            .I(N__38323));
    LocalMux I__8236 (
            .O(N__38329),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__8235 (
            .O(N__38326),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__8234 (
            .O(N__38323),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__8233 (
            .O(N__38316),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__8232 (
            .O(N__38313),
            .I(N__38308));
    InMux I__8231 (
            .O(N__38312),
            .I(N__38305));
    InMux I__8230 (
            .O(N__38311),
            .I(N__38302));
    InMux I__8229 (
            .O(N__38308),
            .I(N__38299));
    LocalMux I__8228 (
            .O(N__38305),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__8227 (
            .O(N__38302),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__8226 (
            .O(N__38299),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__8225 (
            .O(N__38292),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__8224 (
            .O(N__38289),
            .I(N__38286));
    LocalMux I__8223 (
            .O(N__38286),
            .I(N__38283));
    Span4Mux_v I__8222 (
            .O(N__38283),
            .I(N__38278));
    InMux I__8221 (
            .O(N__38282),
            .I(N__38275));
    InMux I__8220 (
            .O(N__38281),
            .I(N__38272));
    Odrv4 I__8219 (
            .O(N__38278),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__8218 (
            .O(N__38275),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__8217 (
            .O(N__38272),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__8216 (
            .O(N__38265),
            .I(bfn_15_19_0_));
    InMux I__8215 (
            .O(N__38262),
            .I(N__38259));
    LocalMux I__8214 (
            .O(N__38259),
            .I(N__38256));
    Span4Mux_v I__8213 (
            .O(N__38256),
            .I(N__38251));
    InMux I__8212 (
            .O(N__38255),
            .I(N__38248));
    InMux I__8211 (
            .O(N__38254),
            .I(N__38245));
    Odrv4 I__8210 (
            .O(N__38251),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__8209 (
            .O(N__38248),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__8208 (
            .O(N__38245),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__8207 (
            .O(N__38238),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CascadeMux I__8206 (
            .O(N__38235),
            .I(N__38230));
    InMux I__8205 (
            .O(N__38234),
            .I(N__38227));
    InMux I__8204 (
            .O(N__38233),
            .I(N__38224));
    InMux I__8203 (
            .O(N__38230),
            .I(N__38221));
    LocalMux I__8202 (
            .O(N__38227),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__8201 (
            .O(N__38224),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__8200 (
            .O(N__38221),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__8199 (
            .O(N__38214),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    CascadeMux I__8198 (
            .O(N__38211),
            .I(N__38206));
    InMux I__8197 (
            .O(N__38210),
            .I(N__38203));
    InMux I__8196 (
            .O(N__38209),
            .I(N__38200));
    InMux I__8195 (
            .O(N__38206),
            .I(N__38197));
    LocalMux I__8194 (
            .O(N__38203),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__8193 (
            .O(N__38200),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__8192 (
            .O(N__38197),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__8191 (
            .O(N__38190),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    CascadeMux I__8190 (
            .O(N__38187),
            .I(N__38182));
    InMux I__8189 (
            .O(N__38186),
            .I(N__38179));
    InMux I__8188 (
            .O(N__38185),
            .I(N__38176));
    InMux I__8187 (
            .O(N__38182),
            .I(N__38173));
    LocalMux I__8186 (
            .O(N__38179),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__8185 (
            .O(N__38176),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__8184 (
            .O(N__38173),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__8183 (
            .O(N__38166),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__8182 (
            .O(N__38163),
            .I(N__38158));
    InMux I__8181 (
            .O(N__38162),
            .I(N__38155));
    InMux I__8180 (
            .O(N__38161),
            .I(N__38152));
    InMux I__8179 (
            .O(N__38158),
            .I(N__38149));
    LocalMux I__8178 (
            .O(N__38155),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__8177 (
            .O(N__38152),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__8176 (
            .O(N__38149),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__8175 (
            .O(N__38142),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    CascadeMux I__8174 (
            .O(N__38139),
            .I(N__38134));
    InMux I__8173 (
            .O(N__38138),
            .I(N__38131));
    InMux I__8172 (
            .O(N__38137),
            .I(N__38128));
    InMux I__8171 (
            .O(N__38134),
            .I(N__38125));
    LocalMux I__8170 (
            .O(N__38131),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__8169 (
            .O(N__38128),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__8168 (
            .O(N__38125),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__8167 (
            .O(N__38118),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__8166 (
            .O(N__38115),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    InMux I__8165 (
            .O(N__38112),
            .I(N__38109));
    LocalMux I__8164 (
            .O(N__38109),
            .I(N__38106));
    Odrv4 I__8163 (
            .O(N__38106),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ));
    InMux I__8162 (
            .O(N__38103),
            .I(N__38100));
    LocalMux I__8161 (
            .O(N__38100),
            .I(N__38097));
    Odrv4 I__8160 (
            .O(N__38097),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ));
    InMux I__8159 (
            .O(N__38094),
            .I(N__38091));
    LocalMux I__8158 (
            .O(N__38091),
            .I(N__38088));
    Odrv4 I__8157 (
            .O(N__38088),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ));
    InMux I__8156 (
            .O(N__38085),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__8155 (
            .O(N__38082),
            .I(N__38079));
    LocalMux I__8154 (
            .O(N__38079),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ));
    InMux I__8153 (
            .O(N__38076),
            .I(N__38072));
    CascadeMux I__8152 (
            .O(N__38075),
            .I(N__38069));
    LocalMux I__8151 (
            .O(N__38072),
            .I(N__38066));
    InMux I__8150 (
            .O(N__38069),
            .I(N__38063));
    Span4Mux_v I__8149 (
            .O(N__38066),
            .I(N__38057));
    LocalMux I__8148 (
            .O(N__38063),
            .I(N__38057));
    InMux I__8147 (
            .O(N__38062),
            .I(N__38053));
    Span4Mux_h I__8146 (
            .O(N__38057),
            .I(N__38050));
    InMux I__8145 (
            .O(N__38056),
            .I(N__38047));
    LocalMux I__8144 (
            .O(N__38053),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    Odrv4 I__8143 (
            .O(N__38050),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    LocalMux I__8142 (
            .O(N__38047),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    InMux I__8141 (
            .O(N__38040),
            .I(N__38037));
    LocalMux I__8140 (
            .O(N__38037),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ));
    InMux I__8139 (
            .O(N__38034),
            .I(N__38031));
    LocalMux I__8138 (
            .O(N__38031),
            .I(N__38028));
    Odrv12 I__8137 (
            .O(N__38028),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ));
    InMux I__8136 (
            .O(N__38025),
            .I(N__38022));
    LocalMux I__8135 (
            .O(N__38022),
            .I(N__38019));
    Odrv4 I__8134 (
            .O(N__38019),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ));
    InMux I__8133 (
            .O(N__38016),
            .I(N__38013));
    LocalMux I__8132 (
            .O(N__38013),
            .I(N__38010));
    Odrv4 I__8131 (
            .O(N__38010),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ));
    InMux I__8130 (
            .O(N__38007),
            .I(N__38004));
    LocalMux I__8129 (
            .O(N__38004),
            .I(N__38001));
    Odrv4 I__8128 (
            .O(N__38001),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ));
    InMux I__8127 (
            .O(N__37998),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__8126 (
            .O(N__37995),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__8125 (
            .O(N__37992),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__8124 (
            .O(N__37989),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__8123 (
            .O(N__37986),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__8122 (
            .O(N__37983),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__8121 (
            .O(N__37980),
            .I(N__37977));
    LocalMux I__8120 (
            .O(N__37977),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__8119 (
            .O(N__37974),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__8118 (
            .O(N__37971),
            .I(bfn_15_15_0_));
    InMux I__8117 (
            .O(N__37968),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__8116 (
            .O(N__37965),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__8115 (
            .O(N__37962),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__8114 (
            .O(N__37959),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__8113 (
            .O(N__37956),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__8112 (
            .O(N__37953),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__8111 (
            .O(N__37950),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__8110 (
            .O(N__37947),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__8109 (
            .O(N__37944),
            .I(bfn_15_14_0_));
    InMux I__8108 (
            .O(N__37941),
            .I(N__37937));
    CascadeMux I__8107 (
            .O(N__37940),
            .I(N__37933));
    LocalMux I__8106 (
            .O(N__37937),
            .I(N__37929));
    InMux I__8105 (
            .O(N__37936),
            .I(N__37925));
    InMux I__8104 (
            .O(N__37933),
            .I(N__37922));
    CascadeMux I__8103 (
            .O(N__37932),
            .I(N__37919));
    Span4Mux_h I__8102 (
            .O(N__37929),
            .I(N__37916));
    InMux I__8101 (
            .O(N__37928),
            .I(N__37913));
    LocalMux I__8100 (
            .O(N__37925),
            .I(N__37910));
    LocalMux I__8099 (
            .O(N__37922),
            .I(N__37907));
    InMux I__8098 (
            .O(N__37919),
            .I(N__37904));
    Span4Mux_v I__8097 (
            .O(N__37916),
            .I(N__37899));
    LocalMux I__8096 (
            .O(N__37913),
            .I(N__37899));
    Span4Mux_h I__8095 (
            .O(N__37910),
            .I(N__37894));
    Span4Mux_h I__8094 (
            .O(N__37907),
            .I(N__37894));
    LocalMux I__8093 (
            .O(N__37904),
            .I(measured_delay_hc_8));
    Odrv4 I__8092 (
            .O(N__37899),
            .I(measured_delay_hc_8));
    Odrv4 I__8091 (
            .O(N__37894),
            .I(measured_delay_hc_8));
    InMux I__8090 (
            .O(N__37887),
            .I(N__37876));
    InMux I__8089 (
            .O(N__37886),
            .I(N__37876));
    InMux I__8088 (
            .O(N__37885),
            .I(N__37871));
    InMux I__8087 (
            .O(N__37884),
            .I(N__37871));
    CascadeMux I__8086 (
            .O(N__37883),
            .I(N__37866));
    InMux I__8085 (
            .O(N__37882),
            .I(N__37862));
    InMux I__8084 (
            .O(N__37881),
            .I(N__37859));
    LocalMux I__8083 (
            .O(N__37876),
            .I(N__37856));
    LocalMux I__8082 (
            .O(N__37871),
            .I(N__37853));
    CascadeMux I__8081 (
            .O(N__37870),
            .I(N__37849));
    CascadeMux I__8080 (
            .O(N__37869),
            .I(N__37845));
    InMux I__8079 (
            .O(N__37866),
            .I(N__37836));
    InMux I__8078 (
            .O(N__37865),
            .I(N__37836));
    LocalMux I__8077 (
            .O(N__37862),
            .I(N__37833));
    LocalMux I__8076 (
            .O(N__37859),
            .I(N__37830));
    Span4Mux_h I__8075 (
            .O(N__37856),
            .I(N__37827));
    Span4Mux_h I__8074 (
            .O(N__37853),
            .I(N__37824));
    InMux I__8073 (
            .O(N__37852),
            .I(N__37821));
    InMux I__8072 (
            .O(N__37849),
            .I(N__37818));
    InMux I__8071 (
            .O(N__37848),
            .I(N__37815));
    InMux I__8070 (
            .O(N__37845),
            .I(N__37810));
    InMux I__8069 (
            .O(N__37844),
            .I(N__37810));
    InMux I__8068 (
            .O(N__37843),
            .I(N__37805));
    InMux I__8067 (
            .O(N__37842),
            .I(N__37805));
    CascadeMux I__8066 (
            .O(N__37841),
            .I(N__37802));
    LocalMux I__8065 (
            .O(N__37836),
            .I(N__37795));
    Span4Mux_h I__8064 (
            .O(N__37833),
            .I(N__37795));
    Span4Mux_v I__8063 (
            .O(N__37830),
            .I(N__37795));
    Span4Mux_h I__8062 (
            .O(N__37827),
            .I(N__37790));
    Span4Mux_v I__8061 (
            .O(N__37824),
            .I(N__37790));
    LocalMux I__8060 (
            .O(N__37821),
            .I(N__37785));
    LocalMux I__8059 (
            .O(N__37818),
            .I(N__37785));
    LocalMux I__8058 (
            .O(N__37815),
            .I(N__37782));
    LocalMux I__8057 (
            .O(N__37810),
            .I(N__37777));
    LocalMux I__8056 (
            .O(N__37805),
            .I(N__37777));
    InMux I__8055 (
            .O(N__37802),
            .I(N__37774));
    Span4Mux_v I__8054 (
            .O(N__37795),
            .I(N__37771));
    Span4Mux_v I__8053 (
            .O(N__37790),
            .I(N__37766));
    Span4Mux_h I__8052 (
            .O(N__37785),
            .I(N__37766));
    Span4Mux_h I__8051 (
            .O(N__37782),
            .I(N__37761));
    Span4Mux_h I__8050 (
            .O(N__37777),
            .I(N__37761));
    LocalMux I__8049 (
            .O(N__37774),
            .I(measured_delay_hc_31));
    Odrv4 I__8048 (
            .O(N__37771),
            .I(measured_delay_hc_31));
    Odrv4 I__8047 (
            .O(N__37766),
            .I(measured_delay_hc_31));
    Odrv4 I__8046 (
            .O(N__37761),
            .I(measured_delay_hc_31));
    InMux I__8045 (
            .O(N__37752),
            .I(N__37748));
    InMux I__8044 (
            .O(N__37751),
            .I(N__37744));
    LocalMux I__8043 (
            .O(N__37748),
            .I(N__37740));
    CascadeMux I__8042 (
            .O(N__37747),
            .I(N__37736));
    LocalMux I__8041 (
            .O(N__37744),
            .I(N__37733));
    InMux I__8040 (
            .O(N__37743),
            .I(N__37730));
    Span4Mux_v I__8039 (
            .O(N__37740),
            .I(N__37727));
    CascadeMux I__8038 (
            .O(N__37739),
            .I(N__37724));
    InMux I__8037 (
            .O(N__37736),
            .I(N__37721));
    Span4Mux_h I__8036 (
            .O(N__37733),
            .I(N__37718));
    LocalMux I__8035 (
            .O(N__37730),
            .I(N__37715));
    Span4Mux_h I__8034 (
            .O(N__37727),
            .I(N__37712));
    InMux I__8033 (
            .O(N__37724),
            .I(N__37709));
    LocalMux I__8032 (
            .O(N__37721),
            .I(measured_delay_hc_5));
    Odrv4 I__8031 (
            .O(N__37718),
            .I(measured_delay_hc_5));
    Odrv12 I__8030 (
            .O(N__37715),
            .I(measured_delay_hc_5));
    Odrv4 I__8029 (
            .O(N__37712),
            .I(measured_delay_hc_5));
    LocalMux I__8028 (
            .O(N__37709),
            .I(measured_delay_hc_5));
    InMux I__8027 (
            .O(N__37698),
            .I(N__37692));
    InMux I__8026 (
            .O(N__37697),
            .I(N__37684));
    InMux I__8025 (
            .O(N__37696),
            .I(N__37684));
    InMux I__8024 (
            .O(N__37695),
            .I(N__37677));
    LocalMux I__8023 (
            .O(N__37692),
            .I(N__37674));
    InMux I__8022 (
            .O(N__37691),
            .I(N__37669));
    InMux I__8021 (
            .O(N__37690),
            .I(N__37669));
    InMux I__8020 (
            .O(N__37689),
            .I(N__37663));
    LocalMux I__8019 (
            .O(N__37684),
            .I(N__37660));
    InMux I__8018 (
            .O(N__37683),
            .I(N__37653));
    InMux I__8017 (
            .O(N__37682),
            .I(N__37653));
    InMux I__8016 (
            .O(N__37681),
            .I(N__37653));
    InMux I__8015 (
            .O(N__37680),
            .I(N__37642));
    LocalMux I__8014 (
            .O(N__37677),
            .I(N__37637));
    Span4Mux_h I__8013 (
            .O(N__37674),
            .I(N__37637));
    LocalMux I__8012 (
            .O(N__37669),
            .I(N__37634));
    InMux I__8011 (
            .O(N__37668),
            .I(N__37627));
    InMux I__8010 (
            .O(N__37667),
            .I(N__37627));
    InMux I__8009 (
            .O(N__37666),
            .I(N__37627));
    LocalMux I__8008 (
            .O(N__37663),
            .I(N__37624));
    Span4Mux_v I__8007 (
            .O(N__37660),
            .I(N__37619));
    LocalMux I__8006 (
            .O(N__37653),
            .I(N__37619));
    InMux I__8005 (
            .O(N__37652),
            .I(N__37614));
    InMux I__8004 (
            .O(N__37651),
            .I(N__37614));
    InMux I__8003 (
            .O(N__37650),
            .I(N__37601));
    InMux I__8002 (
            .O(N__37649),
            .I(N__37601));
    InMux I__8001 (
            .O(N__37648),
            .I(N__37601));
    InMux I__8000 (
            .O(N__37647),
            .I(N__37601));
    InMux I__7999 (
            .O(N__37646),
            .I(N__37601));
    InMux I__7998 (
            .O(N__37645),
            .I(N__37601));
    LocalMux I__7997 (
            .O(N__37642),
            .I(N__37598));
    Span4Mux_v I__7996 (
            .O(N__37637),
            .I(N__37595));
    Span4Mux_h I__7995 (
            .O(N__37634),
            .I(N__37592));
    LocalMux I__7994 (
            .O(N__37627),
            .I(N__37589));
    Span4Mux_v I__7993 (
            .O(N__37624),
            .I(N__37582));
    Span4Mux_h I__7992 (
            .O(N__37619),
            .I(N__37582));
    LocalMux I__7991 (
            .O(N__37614),
            .I(N__37582));
    LocalMux I__7990 (
            .O(N__37601),
            .I(N__37579));
    Odrv12 I__7989 (
            .O(N__37598),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__7988 (
            .O(N__37595),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__7987 (
            .O(N__37592),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv12 I__7986 (
            .O(N__37589),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__7985 (
            .O(N__37582),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv12 I__7984 (
            .O(N__37579),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    CascadeMux I__7983 (
            .O(N__37566),
            .I(N__37563));
    InMux I__7982 (
            .O(N__37563),
            .I(N__37557));
    CascadeMux I__7981 (
            .O(N__37562),
            .I(N__37554));
    InMux I__7980 (
            .O(N__37561),
            .I(N__37551));
    CascadeMux I__7979 (
            .O(N__37560),
            .I(N__37547));
    LocalMux I__7978 (
            .O(N__37557),
            .I(N__37544));
    InMux I__7977 (
            .O(N__37554),
            .I(N__37541));
    LocalMux I__7976 (
            .O(N__37551),
            .I(N__37538));
    CascadeMux I__7975 (
            .O(N__37550),
            .I(N__37535));
    InMux I__7974 (
            .O(N__37547),
            .I(N__37532));
    Span4Mux_h I__7973 (
            .O(N__37544),
            .I(N__37527));
    LocalMux I__7972 (
            .O(N__37541),
            .I(N__37527));
    Span4Mux_h I__7971 (
            .O(N__37538),
            .I(N__37524));
    InMux I__7970 (
            .O(N__37535),
            .I(N__37521));
    LocalMux I__7969 (
            .O(N__37532),
            .I(measured_delay_hc_13));
    Odrv4 I__7968 (
            .O(N__37527),
            .I(measured_delay_hc_13));
    Odrv4 I__7967 (
            .O(N__37524),
            .I(measured_delay_hc_13));
    LocalMux I__7966 (
            .O(N__37521),
            .I(measured_delay_hc_13));
    InMux I__7965 (
            .O(N__37512),
            .I(N__37499));
    InMux I__7964 (
            .O(N__37511),
            .I(N__37499));
    InMux I__7963 (
            .O(N__37510),
            .I(N__37499));
    InMux I__7962 (
            .O(N__37509),
            .I(N__37499));
    InMux I__7961 (
            .O(N__37508),
            .I(N__37496));
    LocalMux I__7960 (
            .O(N__37499),
            .I(N__37492));
    LocalMux I__7959 (
            .O(N__37496),
            .I(N__37489));
    InMux I__7958 (
            .O(N__37495),
            .I(N__37486));
    Span4Mux_v I__7957 (
            .O(N__37492),
            .I(N__37478));
    Span4Mux_h I__7956 (
            .O(N__37489),
            .I(N__37478));
    LocalMux I__7955 (
            .O(N__37486),
            .I(N__37478));
    InMux I__7954 (
            .O(N__37485),
            .I(N__37475));
    Span4Mux_h I__7953 (
            .O(N__37478),
            .I(N__37464));
    LocalMux I__7952 (
            .O(N__37475),
            .I(N__37464));
    InMux I__7951 (
            .O(N__37474),
            .I(N__37461));
    InMux I__7950 (
            .O(N__37473),
            .I(N__37452));
    InMux I__7949 (
            .O(N__37472),
            .I(N__37452));
    InMux I__7948 (
            .O(N__37471),
            .I(N__37452));
    InMux I__7947 (
            .O(N__37470),
            .I(N__37452));
    InMux I__7946 (
            .O(N__37469),
            .I(N__37449));
    Odrv4 I__7945 (
            .O(N__37464),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0 ));
    LocalMux I__7944 (
            .O(N__37461),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0 ));
    LocalMux I__7943 (
            .O(N__37452),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0 ));
    LocalMux I__7942 (
            .O(N__37449),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0 ));
    CascadeMux I__7941 (
            .O(N__37440),
            .I(N__37433));
    CascadeMux I__7940 (
            .O(N__37439),
            .I(N__37430));
    CascadeMux I__7939 (
            .O(N__37438),
            .I(N__37425));
    CascadeMux I__7938 (
            .O(N__37437),
            .I(N__37418));
    CascadeMux I__7937 (
            .O(N__37436),
            .I(N__37413));
    InMux I__7936 (
            .O(N__37433),
            .I(N__37402));
    InMux I__7935 (
            .O(N__37430),
            .I(N__37402));
    InMux I__7934 (
            .O(N__37429),
            .I(N__37402));
    InMux I__7933 (
            .O(N__37428),
            .I(N__37389));
    InMux I__7932 (
            .O(N__37425),
            .I(N__37389));
    InMux I__7931 (
            .O(N__37424),
            .I(N__37389));
    InMux I__7930 (
            .O(N__37423),
            .I(N__37389));
    InMux I__7929 (
            .O(N__37422),
            .I(N__37389));
    InMux I__7928 (
            .O(N__37421),
            .I(N__37389));
    InMux I__7927 (
            .O(N__37418),
            .I(N__37378));
    InMux I__7926 (
            .O(N__37417),
            .I(N__37378));
    InMux I__7925 (
            .O(N__37416),
            .I(N__37378));
    InMux I__7924 (
            .O(N__37413),
            .I(N__37378));
    InMux I__7923 (
            .O(N__37412),
            .I(N__37378));
    InMux I__7922 (
            .O(N__37411),
            .I(N__37375));
    InMux I__7921 (
            .O(N__37410),
            .I(N__37368));
    CascadeMux I__7920 (
            .O(N__37409),
            .I(N__37362));
    LocalMux I__7919 (
            .O(N__37402),
            .I(N__37358));
    LocalMux I__7918 (
            .O(N__37389),
            .I(N__37353));
    LocalMux I__7917 (
            .O(N__37378),
            .I(N__37353));
    LocalMux I__7916 (
            .O(N__37375),
            .I(N__37350));
    InMux I__7915 (
            .O(N__37374),
            .I(N__37346));
    InMux I__7914 (
            .O(N__37373),
            .I(N__37339));
    InMux I__7913 (
            .O(N__37372),
            .I(N__37339));
    InMux I__7912 (
            .O(N__37371),
            .I(N__37339));
    LocalMux I__7911 (
            .O(N__37368),
            .I(N__37336));
    CascadeMux I__7910 (
            .O(N__37367),
            .I(N__37333));
    CascadeMux I__7909 (
            .O(N__37366),
            .I(N__37330));
    CascadeMux I__7908 (
            .O(N__37365),
            .I(N__37325));
    InMux I__7907 (
            .O(N__37362),
            .I(N__37318));
    InMux I__7906 (
            .O(N__37361),
            .I(N__37315));
    Span4Mux_v I__7905 (
            .O(N__37358),
            .I(N__37310));
    Span4Mux_v I__7904 (
            .O(N__37353),
            .I(N__37310));
    Span4Mux_h I__7903 (
            .O(N__37350),
            .I(N__37307));
    InMux I__7902 (
            .O(N__37349),
            .I(N__37304));
    LocalMux I__7901 (
            .O(N__37346),
            .I(N__37299));
    LocalMux I__7900 (
            .O(N__37339),
            .I(N__37299));
    Span4Mux_h I__7899 (
            .O(N__37336),
            .I(N__37296));
    InMux I__7898 (
            .O(N__37333),
            .I(N__37293));
    InMux I__7897 (
            .O(N__37330),
            .I(N__37288));
    InMux I__7896 (
            .O(N__37329),
            .I(N__37288));
    InMux I__7895 (
            .O(N__37328),
            .I(N__37275));
    InMux I__7894 (
            .O(N__37325),
            .I(N__37275));
    InMux I__7893 (
            .O(N__37324),
            .I(N__37275));
    InMux I__7892 (
            .O(N__37323),
            .I(N__37275));
    InMux I__7891 (
            .O(N__37322),
            .I(N__37275));
    InMux I__7890 (
            .O(N__37321),
            .I(N__37275));
    LocalMux I__7889 (
            .O(N__37318),
            .I(N__37270));
    LocalMux I__7888 (
            .O(N__37315),
            .I(N__37270));
    Span4Mux_h I__7887 (
            .O(N__37310),
            .I(N__37267));
    Span4Mux_h I__7886 (
            .O(N__37307),
            .I(N__37264));
    LocalMux I__7885 (
            .O(N__37304),
            .I(N__37257));
    Span4Mux_h I__7884 (
            .O(N__37299),
            .I(N__37257));
    Span4Mux_h I__7883 (
            .O(N__37296),
            .I(N__37257));
    LocalMux I__7882 (
            .O(N__37293),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__7881 (
            .O(N__37288),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__7880 (
            .O(N__37275),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__7879 (
            .O(N__37270),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__7878 (
            .O(N__37267),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__7877 (
            .O(N__37264),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__7876 (
            .O(N__37257),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__7875 (
            .O(N__37242),
            .I(N__37238));
    CascadeMux I__7874 (
            .O(N__37241),
            .I(N__37235));
    InMux I__7873 (
            .O(N__37238),
            .I(N__37230));
    InMux I__7872 (
            .O(N__37235),
            .I(N__37227));
    InMux I__7871 (
            .O(N__37234),
            .I(N__37224));
    CascadeMux I__7870 (
            .O(N__37233),
            .I(N__37220));
    LocalMux I__7869 (
            .O(N__37230),
            .I(N__37217));
    LocalMux I__7868 (
            .O(N__37227),
            .I(N__37214));
    LocalMux I__7867 (
            .O(N__37224),
            .I(N__37211));
    InMux I__7866 (
            .O(N__37223),
            .I(N__37208));
    InMux I__7865 (
            .O(N__37220),
            .I(N__37205));
    Span4Mux_h I__7864 (
            .O(N__37217),
            .I(N__37196));
    Span4Mux_h I__7863 (
            .O(N__37214),
            .I(N__37196));
    Span4Mux_v I__7862 (
            .O(N__37211),
            .I(N__37196));
    LocalMux I__7861 (
            .O(N__37208),
            .I(N__37196));
    LocalMux I__7860 (
            .O(N__37205),
            .I(measured_delay_hc_7));
    Odrv4 I__7859 (
            .O(N__37196),
            .I(measured_delay_hc_7));
    InMux I__7858 (
            .O(N__37191),
            .I(N__37181));
    InMux I__7857 (
            .O(N__37190),
            .I(N__37181));
    InMux I__7856 (
            .O(N__37189),
            .I(N__37176));
    InMux I__7855 (
            .O(N__37188),
            .I(N__37176));
    InMux I__7854 (
            .O(N__37187),
            .I(N__37173));
    InMux I__7853 (
            .O(N__37186),
            .I(N__37170));
    LocalMux I__7852 (
            .O(N__37181),
            .I(N__37163));
    LocalMux I__7851 (
            .O(N__37176),
            .I(N__37163));
    LocalMux I__7850 (
            .O(N__37173),
            .I(N__37163));
    LocalMux I__7849 (
            .O(N__37170),
            .I(N__37157));
    Span4Mux_v I__7848 (
            .O(N__37163),
            .I(N__37150));
    InMux I__7847 (
            .O(N__37162),
            .I(N__37145));
    InMux I__7846 (
            .O(N__37161),
            .I(N__37145));
    InMux I__7845 (
            .O(N__37160),
            .I(N__37142));
    Span4Mux_v I__7844 (
            .O(N__37157),
            .I(N__37138));
    InMux I__7843 (
            .O(N__37156),
            .I(N__37133));
    InMux I__7842 (
            .O(N__37155),
            .I(N__37133));
    InMux I__7841 (
            .O(N__37154),
            .I(N__37128));
    InMux I__7840 (
            .O(N__37153),
            .I(N__37128));
    Span4Mux_h I__7839 (
            .O(N__37150),
            .I(N__37121));
    LocalMux I__7838 (
            .O(N__37145),
            .I(N__37121));
    LocalMux I__7837 (
            .O(N__37142),
            .I(N__37121));
    InMux I__7836 (
            .O(N__37141),
            .I(N__37118));
    Odrv4 I__7835 (
            .O(N__37138),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0 ));
    LocalMux I__7834 (
            .O(N__37133),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0 ));
    LocalMux I__7833 (
            .O(N__37128),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0 ));
    Odrv4 I__7832 (
            .O(N__37121),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0 ));
    LocalMux I__7831 (
            .O(N__37118),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0 ));
    CEMux I__7830 (
            .O(N__37107),
            .I(N__37103));
    CEMux I__7829 (
            .O(N__37106),
            .I(N__37100));
    LocalMux I__7828 (
            .O(N__37103),
            .I(N__37096));
    LocalMux I__7827 (
            .O(N__37100),
            .I(N__37093));
    CEMux I__7826 (
            .O(N__37099),
            .I(N__37088));
    Span4Mux_v I__7825 (
            .O(N__37096),
            .I(N__37083));
    Span4Mux_v I__7824 (
            .O(N__37093),
            .I(N__37083));
    CEMux I__7823 (
            .O(N__37092),
            .I(N__37080));
    CEMux I__7822 (
            .O(N__37091),
            .I(N__37077));
    LocalMux I__7821 (
            .O(N__37088),
            .I(N__37074));
    Span4Mux_h I__7820 (
            .O(N__37083),
            .I(N__37071));
    LocalMux I__7819 (
            .O(N__37080),
            .I(N__37068));
    LocalMux I__7818 (
            .O(N__37077),
            .I(N__37065));
    Span4Mux_v I__7817 (
            .O(N__37074),
            .I(N__37062));
    Span4Mux_h I__7816 (
            .O(N__37071),
            .I(N__37057));
    Span4Mux_v I__7815 (
            .O(N__37068),
            .I(N__37057));
    Span4Mux_v I__7814 (
            .O(N__37065),
            .I(N__37052));
    Span4Mux_v I__7813 (
            .O(N__37062),
            .I(N__37052));
    Odrv4 I__7812 (
            .O(N__37057),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__7811 (
            .O(N__37052),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__7810 (
            .O(N__37047),
            .I(N__37043));
    InMux I__7809 (
            .O(N__37046),
            .I(N__37039));
    LocalMux I__7808 (
            .O(N__37043),
            .I(N__37033));
    InMux I__7807 (
            .O(N__37042),
            .I(N__37030));
    LocalMux I__7806 (
            .O(N__37039),
            .I(N__37027));
    InMux I__7805 (
            .O(N__37038),
            .I(N__37024));
    InMux I__7804 (
            .O(N__37037),
            .I(N__37021));
    InMux I__7803 (
            .O(N__37036),
            .I(N__37018));
    Span4Mux_h I__7802 (
            .O(N__37033),
            .I(N__37013));
    LocalMux I__7801 (
            .O(N__37030),
            .I(N__37013));
    Span12Mux_s8_v I__7800 (
            .O(N__37027),
            .I(N__37010));
    LocalMux I__7799 (
            .O(N__37024),
            .I(N__37007));
    LocalMux I__7798 (
            .O(N__37021),
            .I(N__37004));
    LocalMux I__7797 (
            .O(N__37018),
            .I(measured_delay_hc_9));
    Odrv4 I__7796 (
            .O(N__37013),
            .I(measured_delay_hc_9));
    Odrv12 I__7795 (
            .O(N__37010),
            .I(measured_delay_hc_9));
    Odrv12 I__7794 (
            .O(N__37007),
            .I(measured_delay_hc_9));
    Odrv4 I__7793 (
            .O(N__37004),
            .I(measured_delay_hc_9));
    CascadeMux I__7792 (
            .O(N__36993),
            .I(N__36989));
    InMux I__7791 (
            .O(N__36992),
            .I(N__36986));
    InMux I__7790 (
            .O(N__36989),
            .I(N__36982));
    LocalMux I__7789 (
            .O(N__36986),
            .I(N__36979));
    InMux I__7788 (
            .O(N__36985),
            .I(N__36975));
    LocalMux I__7787 (
            .O(N__36982),
            .I(N__36972));
    Span4Mux_h I__7786 (
            .O(N__36979),
            .I(N__36969));
    InMux I__7785 (
            .O(N__36978),
            .I(N__36966));
    LocalMux I__7784 (
            .O(N__36975),
            .I(measured_delay_hc_0));
    Odrv12 I__7783 (
            .O(N__36972),
            .I(measured_delay_hc_0));
    Odrv4 I__7782 (
            .O(N__36969),
            .I(measured_delay_hc_0));
    LocalMux I__7781 (
            .O(N__36966),
            .I(measured_delay_hc_0));
    InMux I__7780 (
            .O(N__36957),
            .I(N__36952));
    CascadeMux I__7779 (
            .O(N__36956),
            .I(N__36948));
    CascadeMux I__7778 (
            .O(N__36955),
            .I(N__36945));
    LocalMux I__7777 (
            .O(N__36952),
            .I(N__36942));
    InMux I__7776 (
            .O(N__36951),
            .I(N__36939));
    InMux I__7775 (
            .O(N__36948),
            .I(N__36935));
    InMux I__7774 (
            .O(N__36945),
            .I(N__36932));
    Span4Mux_h I__7773 (
            .O(N__36942),
            .I(N__36927));
    LocalMux I__7772 (
            .O(N__36939),
            .I(N__36927));
    InMux I__7771 (
            .O(N__36938),
            .I(N__36924));
    LocalMux I__7770 (
            .O(N__36935),
            .I(measured_delay_hc_6));
    LocalMux I__7769 (
            .O(N__36932),
            .I(measured_delay_hc_6));
    Odrv4 I__7768 (
            .O(N__36927),
            .I(measured_delay_hc_6));
    LocalMux I__7767 (
            .O(N__36924),
            .I(measured_delay_hc_6));
    InMux I__7766 (
            .O(N__36915),
            .I(N__36910));
    InMux I__7765 (
            .O(N__36914),
            .I(N__36906));
    InMux I__7764 (
            .O(N__36913),
            .I(N__36903));
    LocalMux I__7763 (
            .O(N__36910),
            .I(N__36900));
    InMux I__7762 (
            .O(N__36909),
            .I(N__36896));
    LocalMux I__7761 (
            .O(N__36906),
            .I(N__36893));
    LocalMux I__7760 (
            .O(N__36903),
            .I(N__36888));
    Span4Mux_v I__7759 (
            .O(N__36900),
            .I(N__36888));
    InMux I__7758 (
            .O(N__36899),
            .I(N__36885));
    LocalMux I__7757 (
            .O(N__36896),
            .I(measured_delay_hc_1));
    Odrv12 I__7756 (
            .O(N__36893),
            .I(measured_delay_hc_1));
    Odrv4 I__7755 (
            .O(N__36888),
            .I(measured_delay_hc_1));
    LocalMux I__7754 (
            .O(N__36885),
            .I(measured_delay_hc_1));
    InMux I__7753 (
            .O(N__36876),
            .I(N__36872));
    InMux I__7752 (
            .O(N__36875),
            .I(N__36868));
    LocalMux I__7751 (
            .O(N__36872),
            .I(N__36864));
    InMux I__7750 (
            .O(N__36871),
            .I(N__36861));
    LocalMux I__7749 (
            .O(N__36868),
            .I(N__36858));
    InMux I__7748 (
            .O(N__36867),
            .I(N__36854));
    Span4Mux_v I__7747 (
            .O(N__36864),
            .I(N__36851));
    LocalMux I__7746 (
            .O(N__36861),
            .I(N__36848));
    Span4Mux_v I__7745 (
            .O(N__36858),
            .I(N__36845));
    InMux I__7744 (
            .O(N__36857),
            .I(N__36842));
    LocalMux I__7743 (
            .O(N__36854),
            .I(measured_delay_hc_3));
    Odrv4 I__7742 (
            .O(N__36851),
            .I(measured_delay_hc_3));
    Odrv12 I__7741 (
            .O(N__36848),
            .I(measured_delay_hc_3));
    Odrv4 I__7740 (
            .O(N__36845),
            .I(measured_delay_hc_3));
    LocalMux I__7739 (
            .O(N__36842),
            .I(measured_delay_hc_3));
    InMux I__7738 (
            .O(N__36831),
            .I(N__36828));
    LocalMux I__7737 (
            .O(N__36828),
            .I(N__36821));
    InMux I__7736 (
            .O(N__36827),
            .I(N__36818));
    InMux I__7735 (
            .O(N__36826),
            .I(N__36815));
    InMux I__7734 (
            .O(N__36825),
            .I(N__36812));
    InMux I__7733 (
            .O(N__36824),
            .I(N__36809));
    Span12Mux_s8_v I__7732 (
            .O(N__36821),
            .I(N__36804));
    LocalMux I__7731 (
            .O(N__36818),
            .I(N__36804));
    LocalMux I__7730 (
            .O(N__36815),
            .I(N__36801));
    LocalMux I__7729 (
            .O(N__36812),
            .I(measured_delay_hc_4));
    LocalMux I__7728 (
            .O(N__36809),
            .I(measured_delay_hc_4));
    Odrv12 I__7727 (
            .O(N__36804),
            .I(measured_delay_hc_4));
    Odrv4 I__7726 (
            .O(N__36801),
            .I(measured_delay_hc_4));
    InMux I__7725 (
            .O(N__36792),
            .I(N__36788));
    InMux I__7724 (
            .O(N__36791),
            .I(N__36785));
    LocalMux I__7723 (
            .O(N__36788),
            .I(N__36779));
    LocalMux I__7722 (
            .O(N__36785),
            .I(N__36779));
    InMux I__7721 (
            .O(N__36784),
            .I(N__36776));
    Span4Mux_v I__7720 (
            .O(N__36779),
            .I(N__36769));
    LocalMux I__7719 (
            .O(N__36776),
            .I(N__36769));
    InMux I__7718 (
            .O(N__36775),
            .I(N__36766));
    InMux I__7717 (
            .O(N__36774),
            .I(N__36763));
    Span4Mux_h I__7716 (
            .O(N__36769),
            .I(N__36760));
    LocalMux I__7715 (
            .O(N__36766),
            .I(measured_delay_hc_16));
    LocalMux I__7714 (
            .O(N__36763),
            .I(measured_delay_hc_16));
    Odrv4 I__7713 (
            .O(N__36760),
            .I(measured_delay_hc_16));
    InMux I__7712 (
            .O(N__36753),
            .I(N__36746));
    InMux I__7711 (
            .O(N__36752),
            .I(N__36743));
    InMux I__7710 (
            .O(N__36751),
            .I(N__36740));
    CascadeMux I__7709 (
            .O(N__36750),
            .I(N__36737));
    InMux I__7708 (
            .O(N__36749),
            .I(N__36734));
    LocalMux I__7707 (
            .O(N__36746),
            .I(N__36731));
    LocalMux I__7706 (
            .O(N__36743),
            .I(N__36728));
    LocalMux I__7705 (
            .O(N__36740),
            .I(N__36725));
    InMux I__7704 (
            .O(N__36737),
            .I(N__36722));
    LocalMux I__7703 (
            .O(N__36734),
            .I(N__36719));
    Span4Mux_h I__7702 (
            .O(N__36731),
            .I(N__36716));
    Span4Mux_h I__7701 (
            .O(N__36728),
            .I(N__36711));
    Span4Mux_h I__7700 (
            .O(N__36725),
            .I(N__36711));
    LocalMux I__7699 (
            .O(N__36722),
            .I(measured_delay_hc_14));
    Odrv4 I__7698 (
            .O(N__36719),
            .I(measured_delay_hc_14));
    Odrv4 I__7697 (
            .O(N__36716),
            .I(measured_delay_hc_14));
    Odrv4 I__7696 (
            .O(N__36711),
            .I(measured_delay_hc_14));
    InMux I__7695 (
            .O(N__36702),
            .I(N__36698));
    InMux I__7694 (
            .O(N__36701),
            .I(N__36694));
    LocalMux I__7693 (
            .O(N__36698),
            .I(N__36690));
    InMux I__7692 (
            .O(N__36697),
            .I(N__36687));
    LocalMux I__7691 (
            .O(N__36694),
            .I(N__36684));
    InMux I__7690 (
            .O(N__36693),
            .I(N__36680));
    Span4Mux_h I__7689 (
            .O(N__36690),
            .I(N__36675));
    LocalMux I__7688 (
            .O(N__36687),
            .I(N__36675));
    Span4Mux_v I__7687 (
            .O(N__36684),
            .I(N__36672));
    InMux I__7686 (
            .O(N__36683),
            .I(N__36669));
    LocalMux I__7685 (
            .O(N__36680),
            .I(measured_delay_hc_10));
    Odrv4 I__7684 (
            .O(N__36675),
            .I(measured_delay_hc_10));
    Odrv4 I__7683 (
            .O(N__36672),
            .I(measured_delay_hc_10));
    LocalMux I__7682 (
            .O(N__36669),
            .I(measured_delay_hc_10));
    CascadeMux I__7681 (
            .O(N__36660),
            .I(N__36657));
    InMux I__7680 (
            .O(N__36657),
            .I(N__36652));
    InMux I__7679 (
            .O(N__36656),
            .I(N__36649));
    InMux I__7678 (
            .O(N__36655),
            .I(N__36645));
    LocalMux I__7677 (
            .O(N__36652),
            .I(N__36640));
    LocalMux I__7676 (
            .O(N__36649),
            .I(N__36640));
    CascadeMux I__7675 (
            .O(N__36648),
            .I(N__36637));
    LocalMux I__7674 (
            .O(N__36645),
            .I(N__36634));
    Span4Mux_v I__7673 (
            .O(N__36640),
            .I(N__36631));
    InMux I__7672 (
            .O(N__36637),
            .I(N__36627));
    Span12Mux_h I__7671 (
            .O(N__36634),
            .I(N__36624));
    Span4Mux_h I__7670 (
            .O(N__36631),
            .I(N__36621));
    InMux I__7669 (
            .O(N__36630),
            .I(N__36618));
    LocalMux I__7668 (
            .O(N__36627),
            .I(measured_delay_hc_11));
    Odrv12 I__7667 (
            .O(N__36624),
            .I(measured_delay_hc_11));
    Odrv4 I__7666 (
            .O(N__36621),
            .I(measured_delay_hc_11));
    LocalMux I__7665 (
            .O(N__36618),
            .I(measured_delay_hc_11));
    InMux I__7664 (
            .O(N__36609),
            .I(N__36603));
    CascadeMux I__7663 (
            .O(N__36608),
            .I(N__36600));
    InMux I__7662 (
            .O(N__36607),
            .I(N__36597));
    InMux I__7661 (
            .O(N__36606),
            .I(N__36594));
    LocalMux I__7660 (
            .O(N__36603),
            .I(N__36591));
    InMux I__7659 (
            .O(N__36600),
            .I(N__36587));
    LocalMux I__7658 (
            .O(N__36597),
            .I(N__36584));
    LocalMux I__7657 (
            .O(N__36594),
            .I(N__36581));
    Span4Mux_h I__7656 (
            .O(N__36591),
            .I(N__36578));
    InMux I__7655 (
            .O(N__36590),
            .I(N__36575));
    LocalMux I__7654 (
            .O(N__36587),
            .I(measured_delay_hc_12));
    Odrv4 I__7653 (
            .O(N__36584),
            .I(measured_delay_hc_12));
    Odrv12 I__7652 (
            .O(N__36581),
            .I(measured_delay_hc_12));
    Odrv4 I__7651 (
            .O(N__36578),
            .I(measured_delay_hc_12));
    LocalMux I__7650 (
            .O(N__36575),
            .I(measured_delay_hc_12));
    InMux I__7649 (
            .O(N__36564),
            .I(N__36559));
    InMux I__7648 (
            .O(N__36563),
            .I(N__36555));
    InMux I__7647 (
            .O(N__36562),
            .I(N__36552));
    LocalMux I__7646 (
            .O(N__36559),
            .I(N__36548));
    InMux I__7645 (
            .O(N__36558),
            .I(N__36545));
    LocalMux I__7644 (
            .O(N__36555),
            .I(N__36540));
    LocalMux I__7643 (
            .O(N__36552),
            .I(N__36540));
    CascadeMux I__7642 (
            .O(N__36551),
            .I(N__36537));
    Span4Mux_h I__7641 (
            .O(N__36548),
            .I(N__36532));
    LocalMux I__7640 (
            .O(N__36545),
            .I(N__36532));
    Span4Mux_v I__7639 (
            .O(N__36540),
            .I(N__36529));
    InMux I__7638 (
            .O(N__36537),
            .I(N__36526));
    Span4Mux_v I__7637 (
            .O(N__36532),
            .I(N__36521));
    Span4Mux_h I__7636 (
            .O(N__36529),
            .I(N__36521));
    LocalMux I__7635 (
            .O(N__36526),
            .I(measured_delay_hc_19));
    Odrv4 I__7634 (
            .O(N__36521),
            .I(measured_delay_hc_19));
    CascadeMux I__7633 (
            .O(N__36516),
            .I(N__36513));
    InMux I__7632 (
            .O(N__36513),
            .I(N__36509));
    CascadeMux I__7631 (
            .O(N__36512),
            .I(N__36505));
    LocalMux I__7630 (
            .O(N__36509),
            .I(N__36502));
    InMux I__7629 (
            .O(N__36508),
            .I(N__36497));
    InMux I__7628 (
            .O(N__36505),
            .I(N__36494));
    Span4Mux_h I__7627 (
            .O(N__36502),
            .I(N__36491));
    InMux I__7626 (
            .O(N__36501),
            .I(N__36488));
    InMux I__7625 (
            .O(N__36500),
            .I(N__36485));
    LocalMux I__7624 (
            .O(N__36497),
            .I(N__36480));
    LocalMux I__7623 (
            .O(N__36494),
            .I(N__36480));
    Span4Mux_h I__7622 (
            .O(N__36491),
            .I(N__36477));
    LocalMux I__7621 (
            .O(N__36488),
            .I(measured_delay_hc_17));
    LocalMux I__7620 (
            .O(N__36485),
            .I(measured_delay_hc_17));
    Odrv12 I__7619 (
            .O(N__36480),
            .I(measured_delay_hc_17));
    Odrv4 I__7618 (
            .O(N__36477),
            .I(measured_delay_hc_17));
    InMux I__7617 (
            .O(N__36468),
            .I(N__36465));
    LocalMux I__7616 (
            .O(N__36465),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__7615 (
            .O(N__36462),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__7614 (
            .O(N__36459),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__7613 (
            .O(N__36456),
            .I(N__36449));
    CascadeMux I__7612 (
            .O(N__36455),
            .I(N__36443));
    CascadeMux I__7611 (
            .O(N__36454),
            .I(N__36440));
    InMux I__7610 (
            .O(N__36453),
            .I(N__36416));
    InMux I__7609 (
            .O(N__36452),
            .I(N__36416));
    InMux I__7608 (
            .O(N__36449),
            .I(N__36416));
    InMux I__7607 (
            .O(N__36448),
            .I(N__36416));
    InMux I__7606 (
            .O(N__36447),
            .I(N__36416));
    InMux I__7605 (
            .O(N__36446),
            .I(N__36416));
    InMux I__7604 (
            .O(N__36443),
            .I(N__36405));
    InMux I__7603 (
            .O(N__36440),
            .I(N__36405));
    InMux I__7602 (
            .O(N__36439),
            .I(N__36405));
    InMux I__7601 (
            .O(N__36438),
            .I(N__36405));
    InMux I__7600 (
            .O(N__36437),
            .I(N__36405));
    InMux I__7599 (
            .O(N__36436),
            .I(N__36400));
    InMux I__7598 (
            .O(N__36435),
            .I(N__36400));
    InMux I__7597 (
            .O(N__36434),
            .I(N__36395));
    InMux I__7596 (
            .O(N__36433),
            .I(N__36395));
    InMux I__7595 (
            .O(N__36432),
            .I(N__36392));
    InMux I__7594 (
            .O(N__36431),
            .I(N__36385));
    InMux I__7593 (
            .O(N__36430),
            .I(N__36385));
    InMux I__7592 (
            .O(N__36429),
            .I(N__36385));
    LocalMux I__7591 (
            .O(N__36416),
            .I(N__36376));
    LocalMux I__7590 (
            .O(N__36405),
            .I(N__36376));
    LocalMux I__7589 (
            .O(N__36400),
            .I(N__36376));
    LocalMux I__7588 (
            .O(N__36395),
            .I(N__36376));
    LocalMux I__7587 (
            .O(N__36392),
            .I(N__36369));
    LocalMux I__7586 (
            .O(N__36385),
            .I(N__36369));
    Span4Mux_v I__7585 (
            .O(N__36376),
            .I(N__36369));
    Odrv4 I__7584 (
            .O(N__36369),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    CEMux I__7583 (
            .O(N__36366),
            .I(N__36362));
    CEMux I__7582 (
            .O(N__36365),
            .I(N__36359));
    LocalMux I__7581 (
            .O(N__36362),
            .I(N__36356));
    LocalMux I__7580 (
            .O(N__36359),
            .I(N__36352));
    Span4Mux_v I__7579 (
            .O(N__36356),
            .I(N__36349));
    CEMux I__7578 (
            .O(N__36355),
            .I(N__36344));
    Span4Mux_h I__7577 (
            .O(N__36352),
            .I(N__36341));
    Span4Mux_h I__7576 (
            .O(N__36349),
            .I(N__36338));
    CEMux I__7575 (
            .O(N__36348),
            .I(N__36335));
    CEMux I__7574 (
            .O(N__36347),
            .I(N__36332));
    LocalMux I__7573 (
            .O(N__36344),
            .I(N__36329));
    Odrv4 I__7572 (
            .O(N__36341),
            .I(\delay_measurement_inst.delay_tr_timer.N_337_i ));
    Odrv4 I__7571 (
            .O(N__36338),
            .I(\delay_measurement_inst.delay_tr_timer.N_337_i ));
    LocalMux I__7570 (
            .O(N__36335),
            .I(\delay_measurement_inst.delay_tr_timer.N_337_i ));
    LocalMux I__7569 (
            .O(N__36332),
            .I(\delay_measurement_inst.delay_tr_timer.N_337_i ));
    Odrv4 I__7568 (
            .O(N__36329),
            .I(\delay_measurement_inst.delay_tr_timer.N_337_i ));
    InMux I__7567 (
            .O(N__36318),
            .I(N__36315));
    LocalMux I__7566 (
            .O(N__36315),
            .I(N__36312));
    Odrv4 I__7565 (
            .O(N__36312),
            .I(delay_tr_input_c));
    InMux I__7564 (
            .O(N__36309),
            .I(N__36306));
    LocalMux I__7563 (
            .O(N__36306),
            .I(delay_tr_d1));
    InMux I__7562 (
            .O(N__36303),
            .I(N__36298));
    InMux I__7561 (
            .O(N__36302),
            .I(N__36295));
    InMux I__7560 (
            .O(N__36301),
            .I(N__36292));
    LocalMux I__7559 (
            .O(N__36298),
            .I(N__36288));
    LocalMux I__7558 (
            .O(N__36295),
            .I(N__36285));
    LocalMux I__7557 (
            .O(N__36292),
            .I(N__36282));
    InMux I__7556 (
            .O(N__36291),
            .I(N__36279));
    Span4Mux_v I__7555 (
            .O(N__36288),
            .I(N__36272));
    Span4Mux_h I__7554 (
            .O(N__36285),
            .I(N__36272));
    Span4Mux_v I__7553 (
            .O(N__36282),
            .I(N__36272));
    LocalMux I__7552 (
            .O(N__36279),
            .I(N__36269));
    Sp12to4 I__7551 (
            .O(N__36272),
            .I(N__36264));
    Span12Mux_h I__7550 (
            .O(N__36269),
            .I(N__36264));
    Odrv12 I__7549 (
            .O(N__36264),
            .I(delay_tr_d2));
    InMux I__7548 (
            .O(N__36261),
            .I(N__36258));
    LocalMux I__7547 (
            .O(N__36258),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__7546 (
            .O(N__36255),
            .I(N__36252));
    LocalMux I__7545 (
            .O(N__36252),
            .I(N__36249));
    Odrv4 I__7544 (
            .O(N__36249),
            .I(\phase_controller_inst1.N_228 ));
    CascadeMux I__7543 (
            .O(N__36246),
            .I(N__36231));
    CascadeMux I__7542 (
            .O(N__36245),
            .I(N__36224));
    CascadeMux I__7541 (
            .O(N__36244),
            .I(N__36221));
    CascadeMux I__7540 (
            .O(N__36243),
            .I(N__36218));
    CascadeMux I__7539 (
            .O(N__36242),
            .I(N__36215));
    InMux I__7538 (
            .O(N__36241),
            .I(N__36212));
    CascadeMux I__7537 (
            .O(N__36240),
            .I(N__36209));
    CascadeMux I__7536 (
            .O(N__36239),
            .I(N__36206));
    CascadeMux I__7535 (
            .O(N__36238),
            .I(N__36203));
    CascadeMux I__7534 (
            .O(N__36237),
            .I(N__36194));
    CascadeMux I__7533 (
            .O(N__36236),
            .I(N__36191));
    CascadeMux I__7532 (
            .O(N__36235),
            .I(N__36188));
    CascadeMux I__7531 (
            .O(N__36234),
            .I(N__36185));
    InMux I__7530 (
            .O(N__36231),
            .I(N__36182));
    InMux I__7529 (
            .O(N__36230),
            .I(N__36179));
    InMux I__7528 (
            .O(N__36229),
            .I(N__36163));
    InMux I__7527 (
            .O(N__36228),
            .I(N__36163));
    InMux I__7526 (
            .O(N__36227),
            .I(N__36163));
    InMux I__7525 (
            .O(N__36224),
            .I(N__36163));
    InMux I__7524 (
            .O(N__36221),
            .I(N__36163));
    InMux I__7523 (
            .O(N__36218),
            .I(N__36163));
    InMux I__7522 (
            .O(N__36215),
            .I(N__36163));
    LocalMux I__7521 (
            .O(N__36212),
            .I(N__36160));
    InMux I__7520 (
            .O(N__36209),
            .I(N__36157));
    InMux I__7519 (
            .O(N__36206),
            .I(N__36146));
    InMux I__7518 (
            .O(N__36203),
            .I(N__36146));
    InMux I__7517 (
            .O(N__36202),
            .I(N__36146));
    InMux I__7516 (
            .O(N__36201),
            .I(N__36146));
    InMux I__7515 (
            .O(N__36200),
            .I(N__36146));
    InMux I__7514 (
            .O(N__36199),
            .I(N__36131));
    InMux I__7513 (
            .O(N__36198),
            .I(N__36131));
    InMux I__7512 (
            .O(N__36197),
            .I(N__36131));
    InMux I__7511 (
            .O(N__36194),
            .I(N__36131));
    InMux I__7510 (
            .O(N__36191),
            .I(N__36131));
    InMux I__7509 (
            .O(N__36188),
            .I(N__36131));
    InMux I__7508 (
            .O(N__36185),
            .I(N__36131));
    LocalMux I__7507 (
            .O(N__36182),
            .I(N__36128));
    LocalMux I__7506 (
            .O(N__36179),
            .I(N__36125));
    CascadeMux I__7505 (
            .O(N__36178),
            .I(N__36122));
    LocalMux I__7504 (
            .O(N__36163),
            .I(N__36119));
    Span4Mux_v I__7503 (
            .O(N__36160),
            .I(N__36116));
    LocalMux I__7502 (
            .O(N__36157),
            .I(N__36105));
    LocalMux I__7501 (
            .O(N__36146),
            .I(N__36105));
    LocalMux I__7500 (
            .O(N__36131),
            .I(N__36105));
    Span4Mux_v I__7499 (
            .O(N__36128),
            .I(N__36105));
    Span4Mux_h I__7498 (
            .O(N__36125),
            .I(N__36105));
    InMux I__7497 (
            .O(N__36122),
            .I(N__36102));
    Span4Mux_h I__7496 (
            .O(N__36119),
            .I(N__36099));
    Span4Mux_h I__7495 (
            .O(N__36116),
            .I(N__36096));
    Span4Mux_v I__7494 (
            .O(N__36105),
            .I(N__36093));
    LocalMux I__7493 (
            .O(N__36102),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__7492 (
            .O(N__36099),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__7491 (
            .O(N__36096),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__7490 (
            .O(N__36093),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__7489 (
            .O(N__36084),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__7488 (
            .O(N__36081),
            .I(N__36078));
    LocalMux I__7487 (
            .O(N__36078),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__7486 (
            .O(N__36075),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__7485 (
            .O(N__36072),
            .I(N__36069));
    LocalMux I__7484 (
            .O(N__36069),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__7483 (
            .O(N__36066),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__7482 (
            .O(N__36063),
            .I(N__36060));
    InMux I__7481 (
            .O(N__36060),
            .I(N__36057));
    LocalMux I__7480 (
            .O(N__36057),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__7479 (
            .O(N__36054),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__7478 (
            .O(N__36051),
            .I(N__36048));
    LocalMux I__7477 (
            .O(N__36048),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__7476 (
            .O(N__36045),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__7475 (
            .O(N__36042),
            .I(N__36039));
    LocalMux I__7474 (
            .O(N__36039),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__7473 (
            .O(N__36036),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__7472 (
            .O(N__36033),
            .I(N__36030));
    LocalMux I__7471 (
            .O(N__36030),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__7470 (
            .O(N__36027),
            .I(bfn_14_23_0_));
    CascadeMux I__7469 (
            .O(N__36024),
            .I(N__36021));
    InMux I__7468 (
            .O(N__36021),
            .I(N__36018));
    LocalMux I__7467 (
            .O(N__36018),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__7466 (
            .O(N__36015),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__7465 (
            .O(N__36012),
            .I(N__36009));
    LocalMux I__7464 (
            .O(N__36009),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__7463 (
            .O(N__36006),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__7462 (
            .O(N__36003),
            .I(N__35999));
    CascadeMux I__7461 (
            .O(N__36002),
            .I(N__35996));
    LocalMux I__7460 (
            .O(N__35999),
            .I(N__35993));
    InMux I__7459 (
            .O(N__35996),
            .I(N__35990));
    Span4Mux_v I__7458 (
            .O(N__35993),
            .I(N__35987));
    LocalMux I__7457 (
            .O(N__35990),
            .I(N__35984));
    Odrv4 I__7456 (
            .O(N__35987),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    Odrv4 I__7455 (
            .O(N__35984),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    InMux I__7454 (
            .O(N__35979),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__7453 (
            .O(N__35976),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__7452 (
            .O(N__35973),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__7451 (
            .O(N__35970),
            .I(N__35967));
    LocalMux I__7450 (
            .O(N__35967),
            .I(N__35962));
    InMux I__7449 (
            .O(N__35966),
            .I(N__35959));
    InMux I__7448 (
            .O(N__35965),
            .I(N__35956));
    Span4Mux_h I__7447 (
            .O(N__35962),
            .I(N__35951));
    LocalMux I__7446 (
            .O(N__35959),
            .I(N__35951));
    LocalMux I__7445 (
            .O(N__35956),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    Odrv4 I__7444 (
            .O(N__35951),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__7443 (
            .O(N__35946),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__7442 (
            .O(N__35943),
            .I(N__35939));
    InMux I__7441 (
            .O(N__35942),
            .I(N__35936));
    InMux I__7440 (
            .O(N__35939),
            .I(N__35933));
    LocalMux I__7439 (
            .O(N__35936),
            .I(N__35929));
    LocalMux I__7438 (
            .O(N__35933),
            .I(N__35926));
    InMux I__7437 (
            .O(N__35932),
            .I(N__35923));
    Span4Mux_v I__7436 (
            .O(N__35929),
            .I(N__35920));
    Span4Mux_h I__7435 (
            .O(N__35926),
            .I(N__35917));
    LocalMux I__7434 (
            .O(N__35923),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv4 I__7433 (
            .O(N__35920),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv4 I__7432 (
            .O(N__35917),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__7431 (
            .O(N__35910),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__7430 (
            .O(N__35907),
            .I(N__35901));
    InMux I__7429 (
            .O(N__35906),
            .I(N__35901));
    LocalMux I__7428 (
            .O(N__35901),
            .I(N__35897));
    InMux I__7427 (
            .O(N__35900),
            .I(N__35894));
    Span4Mux_h I__7426 (
            .O(N__35897),
            .I(N__35891));
    LocalMux I__7425 (
            .O(N__35894),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv4 I__7424 (
            .O(N__35891),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    InMux I__7423 (
            .O(N__35886),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__7422 (
            .O(N__35883),
            .I(N__35879));
    InMux I__7421 (
            .O(N__35882),
            .I(N__35873));
    InMux I__7420 (
            .O(N__35879),
            .I(N__35873));
    InMux I__7419 (
            .O(N__35878),
            .I(N__35870));
    LocalMux I__7418 (
            .O(N__35873),
            .I(N__35867));
    LocalMux I__7417 (
            .O(N__35870),
            .I(N__35862));
    Span4Mux_h I__7416 (
            .O(N__35867),
            .I(N__35862));
    Odrv4 I__7415 (
            .O(N__35862),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    InMux I__7414 (
            .O(N__35859),
            .I(bfn_14_22_0_));
    CascadeMux I__7413 (
            .O(N__35856),
            .I(N__35853));
    InMux I__7412 (
            .O(N__35853),
            .I(N__35850));
    LocalMux I__7411 (
            .O(N__35850),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__7410 (
            .O(N__35847),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__7409 (
            .O(N__35844),
            .I(N__35841));
    LocalMux I__7408 (
            .O(N__35841),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__7407 (
            .O(N__35838),
            .I(N__35834));
    InMux I__7406 (
            .O(N__35837),
            .I(N__35831));
    LocalMux I__7405 (
            .O(N__35834),
            .I(N__35826));
    LocalMux I__7404 (
            .O(N__35831),
            .I(N__35826));
    Odrv4 I__7403 (
            .O(N__35826),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__7402 (
            .O(N__35823),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__7401 (
            .O(N__35820),
            .I(N__35814));
    InMux I__7400 (
            .O(N__35819),
            .I(N__35809));
    InMux I__7399 (
            .O(N__35818),
            .I(N__35809));
    InMux I__7398 (
            .O(N__35817),
            .I(N__35806));
    LocalMux I__7397 (
            .O(N__35814),
            .I(N__35803));
    LocalMux I__7396 (
            .O(N__35809),
            .I(N__35798));
    LocalMux I__7395 (
            .O(N__35806),
            .I(N__35798));
    Odrv4 I__7394 (
            .O(N__35803),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    Odrv4 I__7393 (
            .O(N__35798),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    InMux I__7392 (
            .O(N__35793),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__7391 (
            .O(N__35790),
            .I(N__35786));
    InMux I__7390 (
            .O(N__35789),
            .I(N__35783));
    LocalMux I__7389 (
            .O(N__35786),
            .I(N__35780));
    LocalMux I__7388 (
            .O(N__35783),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    Odrv12 I__7387 (
            .O(N__35780),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__7386 (
            .O(N__35775),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__7385 (
            .O(N__35772),
            .I(N__35769));
    InMux I__7384 (
            .O(N__35769),
            .I(N__35765));
    InMux I__7383 (
            .O(N__35768),
            .I(N__35762));
    LocalMux I__7382 (
            .O(N__35765),
            .I(N__35759));
    LocalMux I__7381 (
            .O(N__35762),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    Odrv4 I__7380 (
            .O(N__35759),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__7379 (
            .O(N__35754),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__7378 (
            .O(N__35751),
            .I(N__35746));
    InMux I__7377 (
            .O(N__35750),
            .I(N__35742));
    CascadeMux I__7376 (
            .O(N__35749),
            .I(N__35738));
    InMux I__7375 (
            .O(N__35746),
            .I(N__35735));
    InMux I__7374 (
            .O(N__35745),
            .I(N__35732));
    LocalMux I__7373 (
            .O(N__35742),
            .I(N__35729));
    InMux I__7372 (
            .O(N__35741),
            .I(N__35726));
    InMux I__7371 (
            .O(N__35738),
            .I(N__35723));
    LocalMux I__7370 (
            .O(N__35735),
            .I(N__35718));
    LocalMux I__7369 (
            .O(N__35732),
            .I(N__35718));
    Span4Mux_h I__7368 (
            .O(N__35729),
            .I(N__35713));
    LocalMux I__7367 (
            .O(N__35726),
            .I(N__35713));
    LocalMux I__7366 (
            .O(N__35723),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    Odrv4 I__7365 (
            .O(N__35718),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    Odrv4 I__7364 (
            .O(N__35713),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    InMux I__7363 (
            .O(N__35706),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__7362 (
            .O(N__35703),
            .I(N__35699));
    InMux I__7361 (
            .O(N__35702),
            .I(N__35696));
    LocalMux I__7360 (
            .O(N__35699),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    LocalMux I__7359 (
            .O(N__35696),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__7358 (
            .O(N__35691),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__7357 (
            .O(N__35688),
            .I(N__35684));
    InMux I__7356 (
            .O(N__35687),
            .I(N__35681));
    LocalMux I__7355 (
            .O(N__35684),
            .I(N__35678));
    LocalMux I__7354 (
            .O(N__35681),
            .I(N__35675));
    Odrv4 I__7353 (
            .O(N__35678),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    Odrv4 I__7352 (
            .O(N__35675),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__7351 (
            .O(N__35670),
            .I(bfn_14_21_0_));
    InMux I__7350 (
            .O(N__35667),
            .I(N__35664));
    LocalMux I__7349 (
            .O(N__35664),
            .I(N__35660));
    InMux I__7348 (
            .O(N__35663),
            .I(N__35657));
    Span4Mux_h I__7347 (
            .O(N__35660),
            .I(N__35654));
    LocalMux I__7346 (
            .O(N__35657),
            .I(N__35651));
    Odrv4 I__7345 (
            .O(N__35654),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    Odrv4 I__7344 (
            .O(N__35651),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__7343 (
            .O(N__35646),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__7342 (
            .O(N__35643),
            .I(\delay_measurement_inst.N_333_cascade_ ));
    InMux I__7341 (
            .O(N__35640),
            .I(N__35636));
    InMux I__7340 (
            .O(N__35639),
            .I(N__35633));
    LocalMux I__7339 (
            .O(N__35636),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    LocalMux I__7338 (
            .O(N__35633),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    InMux I__7337 (
            .O(N__35628),
            .I(N__35623));
    InMux I__7336 (
            .O(N__35627),
            .I(N__35620));
    InMux I__7335 (
            .O(N__35626),
            .I(N__35617));
    LocalMux I__7334 (
            .O(N__35623),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    LocalMux I__7333 (
            .O(N__35620),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    LocalMux I__7332 (
            .O(N__35617),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    InMux I__7331 (
            .O(N__35610),
            .I(N__35595));
    InMux I__7330 (
            .O(N__35609),
            .I(N__35595));
    InMux I__7329 (
            .O(N__35608),
            .I(N__35595));
    InMux I__7328 (
            .O(N__35607),
            .I(N__35595));
    InMux I__7327 (
            .O(N__35606),
            .I(N__35595));
    LocalMux I__7326 (
            .O(N__35595),
            .I(\delay_measurement_inst.N_333 ));
    InMux I__7325 (
            .O(N__35592),
            .I(N__35588));
    InMux I__7324 (
            .O(N__35591),
            .I(N__35585));
    LocalMux I__7323 (
            .O(N__35588),
            .I(N__35580));
    LocalMux I__7322 (
            .O(N__35585),
            .I(N__35580));
    Span4Mux_v I__7321 (
            .O(N__35580),
            .I(N__35577));
    Span4Mux_h I__7320 (
            .O(N__35577),
            .I(N__35573));
    InMux I__7319 (
            .O(N__35576),
            .I(N__35570));
    Odrv4 I__7318 (
            .O(N__35573),
            .I(\delay_measurement_inst.N_328 ));
    LocalMux I__7317 (
            .O(N__35570),
            .I(\delay_measurement_inst.N_328 ));
    CascadeMux I__7316 (
            .O(N__35565),
            .I(N__35558));
    CascadeMux I__7315 (
            .O(N__35564),
            .I(N__35554));
    CascadeMux I__7314 (
            .O(N__35563),
            .I(N__35551));
    InMux I__7313 (
            .O(N__35562),
            .I(N__35544));
    InMux I__7312 (
            .O(N__35561),
            .I(N__35544));
    InMux I__7311 (
            .O(N__35558),
            .I(N__35541));
    InMux I__7310 (
            .O(N__35557),
            .I(N__35530));
    InMux I__7309 (
            .O(N__35554),
            .I(N__35530));
    InMux I__7308 (
            .O(N__35551),
            .I(N__35530));
    InMux I__7307 (
            .O(N__35550),
            .I(N__35530));
    InMux I__7306 (
            .O(N__35549),
            .I(N__35530));
    LocalMux I__7305 (
            .O(N__35544),
            .I(N__35527));
    LocalMux I__7304 (
            .O(N__35541),
            .I(N__35522));
    LocalMux I__7303 (
            .O(N__35530),
            .I(N__35522));
    Span4Mux_h I__7302 (
            .O(N__35527),
            .I(N__35519));
    Span4Mux_v I__7301 (
            .O(N__35522),
            .I(N__35516));
    Odrv4 I__7300 (
            .O(N__35519),
            .I(\delay_measurement_inst.N_324 ));
    Odrv4 I__7299 (
            .O(N__35516),
            .I(\delay_measurement_inst.N_324 ));
    CEMux I__7298 (
            .O(N__35511),
            .I(N__35504));
    CEMux I__7297 (
            .O(N__35510),
            .I(N__35501));
    CEMux I__7296 (
            .O(N__35509),
            .I(N__35498));
    CEMux I__7295 (
            .O(N__35508),
            .I(N__35495));
    CEMux I__7294 (
            .O(N__35507),
            .I(N__35492));
    LocalMux I__7293 (
            .O(N__35504),
            .I(N__35489));
    LocalMux I__7292 (
            .O(N__35501),
            .I(N__35486));
    LocalMux I__7291 (
            .O(N__35498),
            .I(N__35483));
    LocalMux I__7290 (
            .O(N__35495),
            .I(N__35480));
    LocalMux I__7289 (
            .O(N__35492),
            .I(N__35477));
    Span4Mux_v I__7288 (
            .O(N__35489),
            .I(N__35472));
    Span4Mux_h I__7287 (
            .O(N__35486),
            .I(N__35472));
    Span4Mux_v I__7286 (
            .O(N__35483),
            .I(N__35467));
    Span4Mux_h I__7285 (
            .O(N__35480),
            .I(N__35467));
    Odrv12 I__7284 (
            .O(N__35477),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    Odrv4 I__7283 (
            .O(N__35472),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    Odrv4 I__7282 (
            .O(N__35467),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    CascadeMux I__7281 (
            .O(N__35460),
            .I(N__35456));
    CascadeMux I__7280 (
            .O(N__35459),
            .I(N__35453));
    InMux I__7279 (
            .O(N__35456),
            .I(N__35449));
    InMux I__7278 (
            .O(N__35453),
            .I(N__35444));
    InMux I__7277 (
            .O(N__35452),
            .I(N__35444));
    LocalMux I__7276 (
            .O(N__35449),
            .I(N__35439));
    LocalMux I__7275 (
            .O(N__35444),
            .I(N__35439));
    Odrv4 I__7274 (
            .O(N__35439),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    InMux I__7273 (
            .O(N__35436),
            .I(N__35432));
    InMux I__7272 (
            .O(N__35435),
            .I(N__35429));
    LocalMux I__7271 (
            .O(N__35432),
            .I(N__35426));
    LocalMux I__7270 (
            .O(N__35429),
            .I(N__35423));
    Odrv12 I__7269 (
            .O(N__35426),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    Odrv4 I__7268 (
            .O(N__35423),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    InMux I__7267 (
            .O(N__35418),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__7266 (
            .O(N__35415),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_ ));
    CascadeMux I__7265 (
            .O(N__35412),
            .I(N__35407));
    InMux I__7264 (
            .O(N__35411),
            .I(N__35403));
    InMux I__7263 (
            .O(N__35410),
            .I(N__35400));
    InMux I__7262 (
            .O(N__35407),
            .I(N__35395));
    InMux I__7261 (
            .O(N__35406),
            .I(N__35395));
    LocalMux I__7260 (
            .O(N__35403),
            .I(N__35392));
    LocalMux I__7259 (
            .O(N__35400),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    LocalMux I__7258 (
            .O(N__35395),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    Odrv4 I__7257 (
            .O(N__35392),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    InMux I__7256 (
            .O(N__35385),
            .I(N__35380));
    InMux I__7255 (
            .O(N__35384),
            .I(N__35377));
    InMux I__7254 (
            .O(N__35383),
            .I(N__35374));
    LocalMux I__7253 (
            .O(N__35380),
            .I(N__35371));
    LocalMux I__7252 (
            .O(N__35377),
            .I(N__35366));
    LocalMux I__7251 (
            .O(N__35374),
            .I(N__35366));
    Span4Mux_h I__7250 (
            .O(N__35371),
            .I(N__35361));
    Span4Mux_v I__7249 (
            .O(N__35366),
            .I(N__35361));
    Span4Mux_h I__7248 (
            .O(N__35361),
            .I(N__35358));
    Sp12to4 I__7247 (
            .O(N__35358),
            .I(N__35355));
    Odrv12 I__7246 (
            .O(N__35355),
            .I(il_min_comp2_D2));
    InMux I__7245 (
            .O(N__35352),
            .I(N__35349));
    LocalMux I__7244 (
            .O(N__35349),
            .I(N__35346));
    Odrv4 I__7243 (
            .O(N__35346),
            .I(\phase_controller_slave.start_timer_tr_0_sqmuxa ));
    InMux I__7242 (
            .O(N__35343),
            .I(N__35340));
    LocalMux I__7241 (
            .O(N__35340),
            .I(N__35336));
    InMux I__7240 (
            .O(N__35339),
            .I(N__35333));
    Span4Mux_h I__7239 (
            .O(N__35336),
            .I(N__35329));
    LocalMux I__7238 (
            .O(N__35333),
            .I(N__35326));
    InMux I__7237 (
            .O(N__35332),
            .I(N__35323));
    Span4Mux_v I__7236 (
            .O(N__35329),
            .I(N__35320));
    Odrv4 I__7235 (
            .O(N__35326),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__7234 (
            .O(N__35323),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__7233 (
            .O(N__35320),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__7232 (
            .O(N__35313),
            .I(N__35309));
    InMux I__7231 (
            .O(N__35312),
            .I(N__35306));
    LocalMux I__7230 (
            .O(N__35309),
            .I(N__35303));
    LocalMux I__7229 (
            .O(N__35306),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv12 I__7228 (
            .O(N__35303),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    CascadeMux I__7227 (
            .O(N__35298),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6_cascade_ ));
    CascadeMux I__7226 (
            .O(N__35295),
            .I(N__35291));
    InMux I__7225 (
            .O(N__35294),
            .I(N__35282));
    InMux I__7224 (
            .O(N__35291),
            .I(N__35279));
    InMux I__7223 (
            .O(N__35290),
            .I(N__35276));
    InMux I__7222 (
            .O(N__35289),
            .I(N__35273));
    InMux I__7221 (
            .O(N__35288),
            .I(N__35270));
    InMux I__7220 (
            .O(N__35287),
            .I(N__35265));
    InMux I__7219 (
            .O(N__35286),
            .I(N__35265));
    InMux I__7218 (
            .O(N__35285),
            .I(N__35262));
    LocalMux I__7217 (
            .O(N__35282),
            .I(N__35259));
    LocalMux I__7216 (
            .O(N__35279),
            .I(N__35256));
    LocalMux I__7215 (
            .O(N__35276),
            .I(N__35251));
    LocalMux I__7214 (
            .O(N__35273),
            .I(N__35251));
    LocalMux I__7213 (
            .O(N__35270),
            .I(\delay_measurement_inst.N_358 ));
    LocalMux I__7212 (
            .O(N__35265),
            .I(\delay_measurement_inst.N_358 ));
    LocalMux I__7211 (
            .O(N__35262),
            .I(\delay_measurement_inst.N_358 ));
    Odrv4 I__7210 (
            .O(N__35259),
            .I(\delay_measurement_inst.N_358 ));
    Odrv12 I__7209 (
            .O(N__35256),
            .I(\delay_measurement_inst.N_358 ));
    Odrv4 I__7208 (
            .O(N__35251),
            .I(\delay_measurement_inst.N_358 ));
    InMux I__7207 (
            .O(N__35238),
            .I(N__35232));
    InMux I__7206 (
            .O(N__35237),
            .I(N__35232));
    LocalMux I__7205 (
            .O(N__35232),
            .I(\delay_measurement_inst.delay_tr_timer.N_331 ));
    CascadeMux I__7204 (
            .O(N__35229),
            .I(\delay_measurement_inst.delay_tr_timer.N_331_cascade_ ));
    CascadeMux I__7203 (
            .O(N__35226),
            .I(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_ ));
    CascadeMux I__7202 (
            .O(N__35223),
            .I(N__35219));
    InMux I__7201 (
            .O(N__35222),
            .I(N__35211));
    InMux I__7200 (
            .O(N__35219),
            .I(N__35211));
    InMux I__7199 (
            .O(N__35218),
            .I(N__35211));
    LocalMux I__7198 (
            .O(N__35211),
            .I(\phase_controller_slave.tr_time_passed ));
    InMux I__7197 (
            .O(N__35208),
            .I(N__35202));
    InMux I__7196 (
            .O(N__35207),
            .I(N__35202));
    LocalMux I__7195 (
            .O(N__35202),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    InMux I__7194 (
            .O(N__35199),
            .I(N__35194));
    InMux I__7193 (
            .O(N__35198),
            .I(N__35189));
    InMux I__7192 (
            .O(N__35197),
            .I(N__35189));
    LocalMux I__7191 (
            .O(N__35194),
            .I(N__35186));
    LocalMux I__7190 (
            .O(N__35189),
            .I(N__35183));
    Span4Mux_v I__7189 (
            .O(N__35186),
            .I(N__35178));
    Span4Mux_v I__7188 (
            .O(N__35183),
            .I(N__35178));
    Span4Mux_v I__7187 (
            .O(N__35178),
            .I(N__35175));
    Odrv4 I__7186 (
            .O(N__35175),
            .I(il_max_comp2_D2));
    InMux I__7185 (
            .O(N__35172),
            .I(N__35169));
    LocalMux I__7184 (
            .O(N__35169),
            .I(\phase_controller_slave.N_211 ));
    CascadeMux I__7183 (
            .O(N__35166),
            .I(N__35162));
    CascadeMux I__7182 (
            .O(N__35165),
            .I(N__35158));
    InMux I__7181 (
            .O(N__35162),
            .I(N__35151));
    InMux I__7180 (
            .O(N__35161),
            .I(N__35151));
    InMux I__7179 (
            .O(N__35158),
            .I(N__35148));
    InMux I__7178 (
            .O(N__35157),
            .I(N__35143));
    InMux I__7177 (
            .O(N__35156),
            .I(N__35143));
    LocalMux I__7176 (
            .O(N__35151),
            .I(N__35140));
    LocalMux I__7175 (
            .O(N__35148),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__7174 (
            .O(N__35143),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    Odrv4 I__7173 (
            .O(N__35140),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    InMux I__7172 (
            .O(N__35133),
            .I(N__35129));
    InMux I__7171 (
            .O(N__35132),
            .I(N__35126));
    LocalMux I__7170 (
            .O(N__35129),
            .I(N__35123));
    LocalMux I__7169 (
            .O(N__35126),
            .I(N__35120));
    Span4Mux_v I__7168 (
            .O(N__35123),
            .I(N__35114));
    Span4Mux_h I__7167 (
            .O(N__35120),
            .I(N__35114));
    InMux I__7166 (
            .O(N__35119),
            .I(N__35111));
    Odrv4 I__7165 (
            .O(N__35114),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__7164 (
            .O(N__35111),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    InMux I__7163 (
            .O(N__35106),
            .I(N__35103));
    LocalMux I__7162 (
            .O(N__35103),
            .I(N__35098));
    InMux I__7161 (
            .O(N__35102),
            .I(N__35095));
    InMux I__7160 (
            .O(N__35101),
            .I(N__35092));
    Span4Mux_v I__7159 (
            .O(N__35098),
            .I(N__35089));
    LocalMux I__7158 (
            .O(N__35095),
            .I(N__35084));
    LocalMux I__7157 (
            .O(N__35092),
            .I(N__35084));
    Span4Mux_h I__7156 (
            .O(N__35089),
            .I(N__35081));
    Span4Mux_v I__7155 (
            .O(N__35084),
            .I(N__35078));
    Odrv4 I__7154 (
            .O(N__35081),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    Odrv4 I__7153 (
            .O(N__35078),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    InMux I__7152 (
            .O(N__35073),
            .I(N__35069));
    InMux I__7151 (
            .O(N__35072),
            .I(N__35066));
    LocalMux I__7150 (
            .O(N__35069),
            .I(N__35060));
    LocalMux I__7149 (
            .O(N__35066),
            .I(N__35060));
    InMux I__7148 (
            .O(N__35065),
            .I(N__35056));
    Span4Mux_s3_v I__7147 (
            .O(N__35060),
            .I(N__35051));
    CascadeMux I__7146 (
            .O(N__35059),
            .I(N__35048));
    LocalMux I__7145 (
            .O(N__35056),
            .I(N__35044));
    InMux I__7144 (
            .O(N__35055),
            .I(N__35041));
    InMux I__7143 (
            .O(N__35054),
            .I(N__35038));
    Span4Mux_h I__7142 (
            .O(N__35051),
            .I(N__35034));
    InMux I__7141 (
            .O(N__35048),
            .I(N__35031));
    InMux I__7140 (
            .O(N__35047),
            .I(N__35028));
    Span4Mux_v I__7139 (
            .O(N__35044),
            .I(N__35023));
    LocalMux I__7138 (
            .O(N__35041),
            .I(N__35023));
    LocalMux I__7137 (
            .O(N__35038),
            .I(N__35020));
    InMux I__7136 (
            .O(N__35037),
            .I(N__35017));
    Sp12to4 I__7135 (
            .O(N__35034),
            .I(N__35014));
    LocalMux I__7134 (
            .O(N__35031),
            .I(N__35009));
    LocalMux I__7133 (
            .O(N__35028),
            .I(N__35009));
    Span4Mux_v I__7132 (
            .O(N__35023),
            .I(N__35002));
    Span4Mux_v I__7131 (
            .O(N__35020),
            .I(N__35002));
    LocalMux I__7130 (
            .O(N__35017),
            .I(N__35002));
    Span12Mux_v I__7129 (
            .O(N__35014),
            .I(N__34999));
    Span4Mux_v I__7128 (
            .O(N__35009),
            .I(N__34996));
    Span4Mux_v I__7127 (
            .O(N__35002),
            .I(N__34993));
    Span12Mux_v I__7126 (
            .O(N__34999),
            .I(N__34988));
    Sp12to4 I__7125 (
            .O(N__34996),
            .I(N__34988));
    Span4Mux_h I__7124 (
            .O(N__34993),
            .I(N__34985));
    Span12Mux_h I__7123 (
            .O(N__34988),
            .I(N__34982));
    Span4Mux_v I__7122 (
            .O(N__34985),
            .I(N__34979));
    Odrv12 I__7121 (
            .O(N__34982),
            .I(start_stop_c));
    Odrv4 I__7120 (
            .O(N__34979),
            .I(start_stop_c));
    InMux I__7119 (
            .O(N__34974),
            .I(N__34964));
    InMux I__7118 (
            .O(N__34973),
            .I(N__34964));
    InMux I__7117 (
            .O(N__34972),
            .I(N__34964));
    InMux I__7116 (
            .O(N__34971),
            .I(N__34961));
    LocalMux I__7115 (
            .O(N__34964),
            .I(N__34958));
    LocalMux I__7114 (
            .O(N__34961),
            .I(N__34955));
    Span4Mux_v I__7113 (
            .O(N__34958),
            .I(N__34952));
    Span4Mux_h I__7112 (
            .O(N__34955),
            .I(N__34949));
    Odrv4 I__7111 (
            .O(N__34952),
            .I(shift_flag_start));
    Odrv4 I__7110 (
            .O(N__34949),
            .I(shift_flag_start));
    InMux I__7109 (
            .O(N__34944),
            .I(N__34938));
    InMux I__7108 (
            .O(N__34943),
            .I(N__34935));
    InMux I__7107 (
            .O(N__34942),
            .I(N__34930));
    InMux I__7106 (
            .O(N__34941),
            .I(N__34930));
    LocalMux I__7105 (
            .O(N__34938),
            .I(N__34927));
    LocalMux I__7104 (
            .O(N__34935),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    LocalMux I__7103 (
            .O(N__34930),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    Odrv4 I__7102 (
            .O(N__34927),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    InMux I__7101 (
            .O(N__34920),
            .I(N__34917));
    LocalMux I__7100 (
            .O(N__34917),
            .I(\phase_controller_slave.N_213 ));
    InMux I__7099 (
            .O(N__34914),
            .I(N__34911));
    LocalMux I__7098 (
            .O(N__34911),
            .I(\phase_controller_slave.start_timer_hc_0_sqmuxa ));
    InMux I__7097 (
            .O(N__34908),
            .I(N__34905));
    LocalMux I__7096 (
            .O(N__34905),
            .I(\phase_controller_slave.N_214 ));
    IoInMux I__7095 (
            .O(N__34902),
            .I(N__34899));
    LocalMux I__7094 (
            .O(N__34899),
            .I(N__34896));
    Span12Mux_s4_v I__7093 (
            .O(N__34896),
            .I(N__34892));
    CascadeMux I__7092 (
            .O(N__34895),
            .I(N__34889));
    Span12Mux_v I__7091 (
            .O(N__34892),
            .I(N__34886));
    InMux I__7090 (
            .O(N__34889),
            .I(N__34883));
    Odrv12 I__7089 (
            .O(N__34886),
            .I(s4_phy_c));
    LocalMux I__7088 (
            .O(N__34883),
            .I(s4_phy_c));
    InMux I__7087 (
            .O(N__34878),
            .I(N__34873));
    InMux I__7086 (
            .O(N__34877),
            .I(N__34870));
    InMux I__7085 (
            .O(N__34876),
            .I(N__34867));
    LocalMux I__7084 (
            .O(N__34873),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    LocalMux I__7083 (
            .O(N__34870),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    LocalMux I__7082 (
            .O(N__34867),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    InMux I__7081 (
            .O(N__34860),
            .I(N__34854));
    InMux I__7080 (
            .O(N__34859),
            .I(N__34851));
    InMux I__7079 (
            .O(N__34858),
            .I(N__34848));
    InMux I__7078 (
            .O(N__34857),
            .I(N__34845));
    LocalMux I__7077 (
            .O(N__34854),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__7076 (
            .O(N__34851),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__7075 (
            .O(N__34848),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__7074 (
            .O(N__34845),
            .I(\phase_controller_slave.hc_time_passed ));
    IoInMux I__7073 (
            .O(N__34836),
            .I(N__34833));
    LocalMux I__7072 (
            .O(N__34833),
            .I(N__34830));
    Span4Mux_s0_v I__7071 (
            .O(N__34830),
            .I(N__34827));
    Sp12to4 I__7070 (
            .O(N__34827),
            .I(N__34824));
    Span12Mux_h I__7069 (
            .O(N__34824),
            .I(N__34820));
    CascadeMux I__7068 (
            .O(N__34823),
            .I(N__34816));
    Span12Mux_v I__7067 (
            .O(N__34820),
            .I(N__34813));
    InMux I__7066 (
            .O(N__34819),
            .I(N__34810));
    InMux I__7065 (
            .O(N__34816),
            .I(N__34807));
    Odrv12 I__7064 (
            .O(N__34813),
            .I(s3_phy_c));
    LocalMux I__7063 (
            .O(N__34810),
            .I(s3_phy_c));
    LocalMux I__7062 (
            .O(N__34807),
            .I(s3_phy_c));
    CascadeMux I__7061 (
            .O(N__34800),
            .I(\phase_controller_slave.N_211_cascade_ ));
    IoInMux I__7060 (
            .O(N__34797),
            .I(N__34794));
    LocalMux I__7059 (
            .O(N__34794),
            .I(N__34790));
    CEMux I__7058 (
            .O(N__34793),
            .I(N__34787));
    IoSpan4Mux I__7057 (
            .O(N__34790),
            .I(N__34782));
    LocalMux I__7056 (
            .O(N__34787),
            .I(N__34778));
    CEMux I__7055 (
            .O(N__34786),
            .I(N__34775));
    CEMux I__7054 (
            .O(N__34785),
            .I(N__34772));
    Span4Mux_s3_v I__7053 (
            .O(N__34782),
            .I(N__34769));
    CEMux I__7052 (
            .O(N__34781),
            .I(N__34766));
    Span4Mux_v I__7051 (
            .O(N__34778),
            .I(N__34761));
    LocalMux I__7050 (
            .O(N__34775),
            .I(N__34761));
    LocalMux I__7049 (
            .O(N__34772),
            .I(N__34758));
    Sp12to4 I__7048 (
            .O(N__34769),
            .I(N__34755));
    LocalMux I__7047 (
            .O(N__34766),
            .I(N__34752));
    Span4Mux_v I__7046 (
            .O(N__34761),
            .I(N__34747));
    Span4Mux_h I__7045 (
            .O(N__34758),
            .I(N__34747));
    Span12Mux_s11_v I__7044 (
            .O(N__34755),
            .I(N__34742));
    Sp12to4 I__7043 (
            .O(N__34752),
            .I(N__34742));
    Span4Mux_v I__7042 (
            .O(N__34747),
            .I(N__34739));
    Odrv12 I__7041 (
            .O(N__34742),
            .I(red_c_i));
    Odrv4 I__7040 (
            .O(N__34739),
            .I(red_c_i));
    InMux I__7039 (
            .O(N__34734),
            .I(N__34731));
    LocalMux I__7038 (
            .O(N__34731),
            .I(N__34726));
    CascadeMux I__7037 (
            .O(N__34730),
            .I(N__34722));
    InMux I__7036 (
            .O(N__34729),
            .I(N__34719));
    Sp12to4 I__7035 (
            .O(N__34726),
            .I(N__34715));
    CascadeMux I__7034 (
            .O(N__34725),
            .I(N__34712));
    InMux I__7033 (
            .O(N__34722),
            .I(N__34709));
    LocalMux I__7032 (
            .O(N__34719),
            .I(N__34706));
    InMux I__7031 (
            .O(N__34718),
            .I(N__34703));
    Span12Mux_v I__7030 (
            .O(N__34715),
            .I(N__34700));
    InMux I__7029 (
            .O(N__34712),
            .I(N__34697));
    LocalMux I__7028 (
            .O(N__34709),
            .I(N__34690));
    Span4Mux_v I__7027 (
            .O(N__34706),
            .I(N__34690));
    LocalMux I__7026 (
            .O(N__34703),
            .I(N__34690));
    Odrv12 I__7025 (
            .O(N__34700),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__7024 (
            .O(N__34697),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__7023 (
            .O(N__34690),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    InMux I__7022 (
            .O(N__34683),
            .I(N__34678));
    InMux I__7021 (
            .O(N__34682),
            .I(N__34675));
    InMux I__7020 (
            .O(N__34681),
            .I(N__34672));
    LocalMux I__7019 (
            .O(N__34678),
            .I(N__34667));
    LocalMux I__7018 (
            .O(N__34675),
            .I(N__34667));
    LocalMux I__7017 (
            .O(N__34672),
            .I(N__34664));
    Span4Mux_v I__7016 (
            .O(N__34667),
            .I(N__34661));
    Odrv12 I__7015 (
            .O(N__34664),
            .I(il_min_comp1_D2));
    Odrv4 I__7014 (
            .O(N__34661),
            .I(il_min_comp1_D2));
    InMux I__7013 (
            .O(N__34656),
            .I(N__34653));
    LocalMux I__7012 (
            .O(N__34653),
            .I(\phase_controller_inst1.N_232 ));
    CascadeMux I__7011 (
            .O(N__34650),
            .I(N__34647));
    InMux I__7010 (
            .O(N__34647),
            .I(N__34644));
    LocalMux I__7009 (
            .O(N__34644),
            .I(N__34641));
    Odrv4 I__7008 (
            .O(N__34641),
            .I(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__7007 (
            .O(N__34638),
            .I(N__34635));
    LocalMux I__7006 (
            .O(N__34635),
            .I(N__34631));
    InMux I__7005 (
            .O(N__34634),
            .I(N__34628));
    Span4Mux_v I__7004 (
            .O(N__34631),
            .I(N__34623));
    LocalMux I__7003 (
            .O(N__34628),
            .I(N__34620));
    InMux I__7002 (
            .O(N__34627),
            .I(N__34617));
    InMux I__7001 (
            .O(N__34626),
            .I(N__34614));
    Odrv4 I__7000 (
            .O(N__34623),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    Odrv4 I__6999 (
            .O(N__34620),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__6998 (
            .O(N__34617),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__6997 (
            .O(N__34614),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    CascadeMux I__6996 (
            .O(N__34605),
            .I(N__34602));
    InMux I__6995 (
            .O(N__34602),
            .I(N__34599));
    LocalMux I__6994 (
            .O(N__34599),
            .I(N__34596));
    Span4Mux_h I__6993 (
            .O(N__34596),
            .I(N__34593));
    Odrv4 I__6992 (
            .O(N__34593),
            .I(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__6991 (
            .O(N__34590),
            .I(N__34586));
    InMux I__6990 (
            .O(N__34589),
            .I(N__34583));
    LocalMux I__6989 (
            .O(N__34586),
            .I(N__34576));
    LocalMux I__6988 (
            .O(N__34583),
            .I(N__34573));
    InMux I__6987 (
            .O(N__34582),
            .I(N__34570));
    InMux I__6986 (
            .O(N__34581),
            .I(N__34563));
    InMux I__6985 (
            .O(N__34580),
            .I(N__34563));
    InMux I__6984 (
            .O(N__34579),
            .I(N__34563));
    Odrv4 I__6983 (
            .O(N__34576),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__6982 (
            .O(N__34573),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__6981 (
            .O(N__34570),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__6980 (
            .O(N__34563),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__6979 (
            .O(N__34554),
            .I(N__34550));
    InMux I__6978 (
            .O(N__34553),
            .I(N__34547));
    LocalMux I__6977 (
            .O(N__34550),
            .I(N__34541));
    LocalMux I__6976 (
            .O(N__34547),
            .I(N__34541));
    InMux I__6975 (
            .O(N__34546),
            .I(N__34538));
    Span4Mux_v I__6974 (
            .O(N__34541),
            .I(N__34533));
    LocalMux I__6973 (
            .O(N__34538),
            .I(N__34533));
    Span4Mux_v I__6972 (
            .O(N__34533),
            .I(N__34530));
    Odrv4 I__6971 (
            .O(N__34530),
            .I(il_max_comp1_D2));
    InMux I__6970 (
            .O(N__34527),
            .I(N__34523));
    CascadeMux I__6969 (
            .O(N__34526),
            .I(N__34518));
    LocalMux I__6968 (
            .O(N__34523),
            .I(N__34515));
    CascadeMux I__6967 (
            .O(N__34522),
            .I(N__34511));
    CascadeMux I__6966 (
            .O(N__34521),
            .I(N__34508));
    InMux I__6965 (
            .O(N__34518),
            .I(N__34505));
    Span4Mux_v I__6964 (
            .O(N__34515),
            .I(N__34502));
    InMux I__6963 (
            .O(N__34514),
            .I(N__34499));
    InMux I__6962 (
            .O(N__34511),
            .I(N__34496));
    InMux I__6961 (
            .O(N__34508),
            .I(N__34493));
    LocalMux I__6960 (
            .O(N__34505),
            .I(N__34490));
    Span4Mux_v I__6959 (
            .O(N__34502),
            .I(N__34487));
    LocalMux I__6958 (
            .O(N__34499),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__6957 (
            .O(N__34496),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__6956 (
            .O(N__34493),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    Odrv12 I__6955 (
            .O(N__34490),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    Odrv4 I__6954 (
            .O(N__34487),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    InMux I__6953 (
            .O(N__34476),
            .I(N__34466));
    InMux I__6952 (
            .O(N__34475),
            .I(N__34466));
    InMux I__6951 (
            .O(N__34474),
            .I(N__34466));
    InMux I__6950 (
            .O(N__34473),
            .I(N__34463));
    LocalMux I__6949 (
            .O(N__34466),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__6948 (
            .O(N__34463),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__6947 (
            .O(N__34458),
            .I(N__34455));
    LocalMux I__6946 (
            .O(N__34455),
            .I(N__34452));
    Span4Mux_v I__6945 (
            .O(N__34452),
            .I(N__34446));
    InMux I__6944 (
            .O(N__34451),
            .I(N__34441));
    InMux I__6943 (
            .O(N__34450),
            .I(N__34441));
    InMux I__6942 (
            .O(N__34449),
            .I(N__34438));
    Odrv4 I__6941 (
            .O(N__34446),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__6940 (
            .O(N__34441),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__6939 (
            .O(N__34438),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    CascadeMux I__6938 (
            .O(N__34431),
            .I(N__34427));
    InMux I__6937 (
            .O(N__34430),
            .I(N__34423));
    InMux I__6936 (
            .O(N__34427),
            .I(N__34419));
    CascadeMux I__6935 (
            .O(N__34426),
            .I(N__34416));
    LocalMux I__6934 (
            .O(N__34423),
            .I(N__34412));
    InMux I__6933 (
            .O(N__34422),
            .I(N__34409));
    LocalMux I__6932 (
            .O(N__34419),
            .I(N__34406));
    InMux I__6931 (
            .O(N__34416),
            .I(N__34403));
    InMux I__6930 (
            .O(N__34415),
            .I(N__34400));
    Span4Mux_h I__6929 (
            .O(N__34412),
            .I(N__34395));
    LocalMux I__6928 (
            .O(N__34409),
            .I(N__34395));
    Span4Mux_v I__6927 (
            .O(N__34406),
            .I(N__34392));
    LocalMux I__6926 (
            .O(N__34403),
            .I(measured_delay_hc_18));
    LocalMux I__6925 (
            .O(N__34400),
            .I(measured_delay_hc_18));
    Odrv4 I__6924 (
            .O(N__34395),
            .I(measured_delay_hc_18));
    Odrv4 I__6923 (
            .O(N__34392),
            .I(measured_delay_hc_18));
    InMux I__6922 (
            .O(N__34383),
            .I(N__34376));
    InMux I__6921 (
            .O(N__34382),
            .I(N__34376));
    InMux I__6920 (
            .O(N__34381),
            .I(N__34373));
    LocalMux I__6919 (
            .O(N__34376),
            .I(N__34370));
    LocalMux I__6918 (
            .O(N__34373),
            .I(N__34365));
    Span4Mux_v I__6917 (
            .O(N__34370),
            .I(N__34362));
    InMux I__6916 (
            .O(N__34369),
            .I(N__34357));
    InMux I__6915 (
            .O(N__34368),
            .I(N__34357));
    Span4Mux_v I__6914 (
            .O(N__34365),
            .I(N__34354));
    Odrv4 I__6913 (
            .O(N__34362),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2 ));
    LocalMux I__6912 (
            .O(N__34357),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2 ));
    Odrv4 I__6911 (
            .O(N__34354),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2 ));
    InMux I__6910 (
            .O(N__34347),
            .I(N__34343));
    InMux I__6909 (
            .O(N__34346),
            .I(N__34340));
    LocalMux I__6908 (
            .O(N__34343),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__6907 (
            .O(N__34340),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__6906 (
            .O(N__34335),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__6905 (
            .O(N__34332),
            .I(N__34329));
    LocalMux I__6904 (
            .O(N__34329),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    CascadeMux I__6903 (
            .O(N__34326),
            .I(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2_cascade_ ));
    InMux I__6902 (
            .O(N__34323),
            .I(N__34320));
    LocalMux I__6901 (
            .O(N__34320),
            .I(N__34317));
    Span4Mux_h I__6900 (
            .O(N__34317),
            .I(N__34314));
    Odrv4 I__6899 (
            .O(N__34314),
            .I(\phase_controller_inst1.stoper_hc.un1_N_4 ));
    InMux I__6898 (
            .O(N__34311),
            .I(N__34308));
    LocalMux I__6897 (
            .O(N__34308),
            .I(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3 ));
    InMux I__6896 (
            .O(N__34305),
            .I(N__34302));
    LocalMux I__6895 (
            .O(N__34302),
            .I(N__34299));
    Span4Mux_h I__6894 (
            .O(N__34299),
            .I(N__34296));
    Odrv4 I__6893 (
            .O(N__34296),
            .I(\phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1 ));
    InMux I__6892 (
            .O(N__34293),
            .I(N__34288));
    InMux I__6891 (
            .O(N__34292),
            .I(N__34284));
    InMux I__6890 (
            .O(N__34291),
            .I(N__34281));
    LocalMux I__6889 (
            .O(N__34288),
            .I(N__34278));
    InMux I__6888 (
            .O(N__34287),
            .I(N__34275));
    LocalMux I__6887 (
            .O(N__34284),
            .I(N__34270));
    LocalMux I__6886 (
            .O(N__34281),
            .I(N__34270));
    Span4Mux_h I__6885 (
            .O(N__34278),
            .I(N__34265));
    LocalMux I__6884 (
            .O(N__34275),
            .I(N__34265));
    Span4Mux_v I__6883 (
            .O(N__34270),
            .I(N__34262));
    Span4Mux_v I__6882 (
            .O(N__34265),
            .I(N__34259));
    Odrv4 I__6881 (
            .O(N__34262),
            .I(delay_hc_d2));
    Odrv4 I__6880 (
            .O(N__34259),
            .I(delay_hc_d2));
    InMux I__6879 (
            .O(N__34254),
            .I(N__34250));
    InMux I__6878 (
            .O(N__34253),
            .I(N__34247));
    LocalMux I__6877 (
            .O(N__34250),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__6876 (
            .O(N__34247),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__6875 (
            .O(N__34242),
            .I(N__34239));
    InMux I__6874 (
            .O(N__34239),
            .I(N__34236));
    LocalMux I__6873 (
            .O(N__34236),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    InMux I__6872 (
            .O(N__34233),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__6871 (
            .O(N__34230),
            .I(N__34226));
    InMux I__6870 (
            .O(N__34229),
            .I(N__34223));
    LocalMux I__6869 (
            .O(N__34226),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__6868 (
            .O(N__34223),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__6867 (
            .O(N__34218),
            .I(N__34215));
    LocalMux I__6866 (
            .O(N__34215),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    InMux I__6865 (
            .O(N__34212),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__6864 (
            .O(N__34209),
            .I(N__34205));
    InMux I__6863 (
            .O(N__34208),
            .I(N__34202));
    LocalMux I__6862 (
            .O(N__34205),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__6861 (
            .O(N__34202),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__6860 (
            .O(N__34197),
            .I(N__34194));
    LocalMux I__6859 (
            .O(N__34194),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__6858 (
            .O(N__34191),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__6857 (
            .O(N__34188),
            .I(N__34184));
    InMux I__6856 (
            .O(N__34187),
            .I(N__34181));
    LocalMux I__6855 (
            .O(N__34184),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__6854 (
            .O(N__34181),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__6853 (
            .O(N__34176),
            .I(N__34173));
    LocalMux I__6852 (
            .O(N__34173),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__6851 (
            .O(N__34170),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__6850 (
            .O(N__34167),
            .I(N__34163));
    InMux I__6849 (
            .O(N__34166),
            .I(N__34160));
    LocalMux I__6848 (
            .O(N__34163),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__6847 (
            .O(N__34160),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__6846 (
            .O(N__34155),
            .I(N__34152));
    InMux I__6845 (
            .O(N__34152),
            .I(N__34149));
    LocalMux I__6844 (
            .O(N__34149),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    InMux I__6843 (
            .O(N__34146),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__6842 (
            .O(N__34143),
            .I(N__34139));
    InMux I__6841 (
            .O(N__34142),
            .I(N__34136));
    LocalMux I__6840 (
            .O(N__34139),
            .I(N__34133));
    LocalMux I__6839 (
            .O(N__34136),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__6838 (
            .O(N__34133),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__6837 (
            .O(N__34128),
            .I(N__34125));
    InMux I__6836 (
            .O(N__34125),
            .I(N__34122));
    LocalMux I__6835 (
            .O(N__34122),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    InMux I__6834 (
            .O(N__34119),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__6833 (
            .O(N__34116),
            .I(N__34112));
    InMux I__6832 (
            .O(N__34115),
            .I(N__34109));
    LocalMux I__6831 (
            .O(N__34112),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__6830 (
            .O(N__34109),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__6829 (
            .O(N__34104),
            .I(N__34101));
    LocalMux I__6828 (
            .O(N__34101),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__6827 (
            .O(N__34098),
            .I(bfn_14_7_0_));
    InMux I__6826 (
            .O(N__34095),
            .I(N__34091));
    InMux I__6825 (
            .O(N__34094),
            .I(N__34088));
    LocalMux I__6824 (
            .O(N__34091),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__6823 (
            .O(N__34088),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__6822 (
            .O(N__34083),
            .I(N__34080));
    LocalMux I__6821 (
            .O(N__34080),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    InMux I__6820 (
            .O(N__34077),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__6819 (
            .O(N__34074),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__6818 (
            .O(N__34071),
            .I(N__34067));
    InMux I__6817 (
            .O(N__34070),
            .I(N__34064));
    LocalMux I__6816 (
            .O(N__34067),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__6815 (
            .O(N__34064),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__6814 (
            .O(N__34059),
            .I(N__34056));
    LocalMux I__6813 (
            .O(N__34056),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__6812 (
            .O(N__34053),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__6811 (
            .O(N__34050),
            .I(N__34046));
    InMux I__6810 (
            .O(N__34049),
            .I(N__34043));
    LocalMux I__6809 (
            .O(N__34046),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__6808 (
            .O(N__34043),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__6807 (
            .O(N__34038),
            .I(N__34035));
    LocalMux I__6806 (
            .O(N__34035),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__6805 (
            .O(N__34032),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__6804 (
            .O(N__34029),
            .I(N__34025));
    InMux I__6803 (
            .O(N__34028),
            .I(N__34022));
    LocalMux I__6802 (
            .O(N__34025),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__6801 (
            .O(N__34022),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__6800 (
            .O(N__34017),
            .I(N__34014));
    InMux I__6799 (
            .O(N__34014),
            .I(N__34011));
    LocalMux I__6798 (
            .O(N__34011),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__6797 (
            .O(N__34008),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__6796 (
            .O(N__34005),
            .I(N__34001));
    InMux I__6795 (
            .O(N__34004),
            .I(N__33998));
    LocalMux I__6794 (
            .O(N__34001),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__6793 (
            .O(N__33998),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__6792 (
            .O(N__33993),
            .I(N__33990));
    LocalMux I__6791 (
            .O(N__33990),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__6790 (
            .O(N__33987),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__6789 (
            .O(N__33984),
            .I(N__33981));
    LocalMux I__6788 (
            .O(N__33981),
            .I(N__33977));
    InMux I__6787 (
            .O(N__33980),
            .I(N__33974));
    Odrv4 I__6786 (
            .O(N__33977),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__6785 (
            .O(N__33974),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__6784 (
            .O(N__33969),
            .I(N__33966));
    LocalMux I__6783 (
            .O(N__33966),
            .I(N__33963));
    Span4Mux_h I__6782 (
            .O(N__33963),
            .I(N__33960));
    Odrv4 I__6781 (
            .O(N__33960),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__6780 (
            .O(N__33957),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__6779 (
            .O(N__33954),
            .I(N__33950));
    InMux I__6778 (
            .O(N__33953),
            .I(N__33947));
    LocalMux I__6777 (
            .O(N__33950),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__6776 (
            .O(N__33947),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__6775 (
            .O(N__33942),
            .I(N__33939));
    LocalMux I__6774 (
            .O(N__33939),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__6773 (
            .O(N__33936),
            .I(bfn_14_6_0_));
    InMux I__6772 (
            .O(N__33933),
            .I(N__33929));
    InMux I__6771 (
            .O(N__33932),
            .I(N__33926));
    LocalMux I__6770 (
            .O(N__33929),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__6769 (
            .O(N__33926),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__6768 (
            .O(N__33921),
            .I(N__33918));
    InMux I__6767 (
            .O(N__33918),
            .I(N__33915));
    LocalMux I__6766 (
            .O(N__33915),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__6765 (
            .O(N__33912),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__6764 (
            .O(N__33909),
            .I(N__33906));
    LocalMux I__6763 (
            .O(N__33906),
            .I(N__33903));
    Span4Mux_v I__6762 (
            .O(N__33903),
            .I(N__33897));
    InMux I__6761 (
            .O(N__33902),
            .I(N__33894));
    InMux I__6760 (
            .O(N__33901),
            .I(N__33889));
    InMux I__6759 (
            .O(N__33900),
            .I(N__33889));
    Odrv4 I__6758 (
            .O(N__33897),
            .I(\delay_measurement_inst.delay_tr_timer.N_296 ));
    LocalMux I__6757 (
            .O(N__33894),
            .I(\delay_measurement_inst.delay_tr_timer.N_296 ));
    LocalMux I__6756 (
            .O(N__33889),
            .I(\delay_measurement_inst.delay_tr_timer.N_296 ));
    CascadeMux I__6755 (
            .O(N__33882),
            .I(\delay_measurement_inst.delay_tr_timer.N_293_cascade_ ));
    InMux I__6754 (
            .O(N__33879),
            .I(N__33876));
    LocalMux I__6753 (
            .O(N__33876),
            .I(N__33873));
    Odrv4 I__6752 (
            .O(N__33873),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ));
    InMux I__6751 (
            .O(N__33870),
            .I(N__33867));
    LocalMux I__6750 (
            .O(N__33867),
            .I(N__33864));
    Odrv12 I__6749 (
            .O(N__33864),
            .I(\delay_measurement_inst.N_307 ));
    IoInMux I__6748 (
            .O(N__33861),
            .I(N__33858));
    LocalMux I__6747 (
            .O(N__33858),
            .I(N__33855));
    Odrv4 I__6746 (
            .O(N__33855),
            .I(s2_phy_c));
    IoInMux I__6745 (
            .O(N__33852),
            .I(N__33849));
    LocalMux I__6744 (
            .O(N__33849),
            .I(N__33846));
    Span4Mux_s3_v I__6743 (
            .O(N__33846),
            .I(N__33843));
    Odrv4 I__6742 (
            .O(N__33843),
            .I(\delay_measurement_inst.delay_hc_timer.N_335_i ));
    InMux I__6741 (
            .O(N__33840),
            .I(N__33837));
    LocalMux I__6740 (
            .O(N__33837),
            .I(N__33834));
    Span4Mux_h I__6739 (
            .O(N__33834),
            .I(N__33831));
    Odrv4 I__6738 (
            .O(N__33831),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    CascadeMux I__6737 (
            .O(N__33828),
            .I(N__33825));
    InMux I__6736 (
            .O(N__33825),
            .I(N__33821));
    InMux I__6735 (
            .O(N__33824),
            .I(N__33817));
    LocalMux I__6734 (
            .O(N__33821),
            .I(N__33814));
    InMux I__6733 (
            .O(N__33820),
            .I(N__33811));
    LocalMux I__6732 (
            .O(N__33817),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__6731 (
            .O(N__33814),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__6730 (
            .O(N__33811),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__6729 (
            .O(N__33804),
            .I(N__33800));
    InMux I__6728 (
            .O(N__33803),
            .I(N__33797));
    LocalMux I__6727 (
            .O(N__33800),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__6726 (
            .O(N__33797),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__6725 (
            .O(N__33792),
            .I(N__33789));
    LocalMux I__6724 (
            .O(N__33789),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__6723 (
            .O(N__33786),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__6722 (
            .O(N__33783),
            .I(N__33780));
    LocalMux I__6721 (
            .O(N__33780),
            .I(N__33777));
    Span4Mux_h I__6720 (
            .O(N__33777),
            .I(N__33774));
    Odrv4 I__6719 (
            .O(N__33774),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ));
    CascadeMux I__6718 (
            .O(N__33771),
            .I(N__33768));
    InMux I__6717 (
            .O(N__33768),
            .I(N__33764));
    InMux I__6716 (
            .O(N__33767),
            .I(N__33761));
    LocalMux I__6715 (
            .O(N__33764),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__6714 (
            .O(N__33761),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__6713 (
            .O(N__33756),
            .I(N__33753));
    InMux I__6712 (
            .O(N__33753),
            .I(N__33750));
    LocalMux I__6711 (
            .O(N__33750),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    CascadeMux I__6710 (
            .O(N__33747),
            .I(\delay_measurement_inst.N_358_cascade_ ));
    InMux I__6709 (
            .O(N__33744),
            .I(N__33739));
    InMux I__6708 (
            .O(N__33743),
            .I(N__33736));
    InMux I__6707 (
            .O(N__33742),
            .I(N__33733));
    LocalMux I__6706 (
            .O(N__33739),
            .I(N__33730));
    LocalMux I__6705 (
            .O(N__33736),
            .I(N__33726));
    LocalMux I__6704 (
            .O(N__33733),
            .I(N__33721));
    Span12Mux_h I__6703 (
            .O(N__33730),
            .I(N__33721));
    InMux I__6702 (
            .O(N__33729),
            .I(N__33718));
    Span12Mux_v I__6701 (
            .O(N__33726),
            .I(N__33715));
    Span12Mux_v I__6700 (
            .O(N__33721),
            .I(N__33712));
    LocalMux I__6699 (
            .O(N__33718),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    Odrv12 I__6698 (
            .O(N__33715),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    Odrv12 I__6697 (
            .O(N__33712),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    InMux I__6696 (
            .O(N__33705),
            .I(N__33702));
    LocalMux I__6695 (
            .O(N__33702),
            .I(N__33698));
    InMux I__6694 (
            .O(N__33701),
            .I(N__33695));
    Span4Mux_h I__6693 (
            .O(N__33698),
            .I(N__33690));
    LocalMux I__6692 (
            .O(N__33695),
            .I(N__33690));
    Span4Mux_v I__6691 (
            .O(N__33690),
            .I(N__33686));
    InMux I__6690 (
            .O(N__33689),
            .I(N__33683));
    Span4Mux_v I__6689 (
            .O(N__33686),
            .I(N__33680));
    LocalMux I__6688 (
            .O(N__33683),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    Odrv4 I__6687 (
            .O(N__33680),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    InMux I__6686 (
            .O(N__33675),
            .I(N__33670));
    InMux I__6685 (
            .O(N__33674),
            .I(N__33667));
    InMux I__6684 (
            .O(N__33673),
            .I(N__33663));
    LocalMux I__6683 (
            .O(N__33670),
            .I(N__33660));
    LocalMux I__6682 (
            .O(N__33667),
            .I(N__33657));
    InMux I__6681 (
            .O(N__33666),
            .I(N__33654));
    LocalMux I__6680 (
            .O(N__33663),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    Odrv12 I__6679 (
            .O(N__33660),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    Odrv4 I__6678 (
            .O(N__33657),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    LocalMux I__6677 (
            .O(N__33654),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    CEMux I__6676 (
            .O(N__33645),
            .I(N__33642));
    LocalMux I__6675 (
            .O(N__33642),
            .I(N__33636));
    CEMux I__6674 (
            .O(N__33641),
            .I(N__33633));
    CEMux I__6673 (
            .O(N__33640),
            .I(N__33630));
    CEMux I__6672 (
            .O(N__33639),
            .I(N__33627));
    Span4Mux_v I__6671 (
            .O(N__33636),
            .I(N__33624));
    LocalMux I__6670 (
            .O(N__33633),
            .I(N__33619));
    LocalMux I__6669 (
            .O(N__33630),
            .I(N__33619));
    LocalMux I__6668 (
            .O(N__33627),
            .I(N__33616));
    Span4Mux_h I__6667 (
            .O(N__33624),
            .I(N__33611));
    Span4Mux_v I__6666 (
            .O(N__33619),
            .I(N__33611));
    Span4Mux_h I__6665 (
            .O(N__33616),
            .I(N__33608));
    Span4Mux_h I__6664 (
            .O(N__33611),
            .I(N__33605));
    Span4Mux_h I__6663 (
            .O(N__33608),
            .I(N__33602));
    Odrv4 I__6662 (
            .O(N__33605),
            .I(\current_shift_inst.timer_phase.N_192_i ));
    Odrv4 I__6661 (
            .O(N__33602),
            .I(\current_shift_inst.timer_phase.N_192_i ));
    InMux I__6660 (
            .O(N__33597),
            .I(N__33594));
    LocalMux I__6659 (
            .O(N__33594),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ));
    InMux I__6658 (
            .O(N__33591),
            .I(N__33588));
    LocalMux I__6657 (
            .O(N__33588),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ));
    InMux I__6656 (
            .O(N__33585),
            .I(N__33579));
    InMux I__6655 (
            .O(N__33584),
            .I(N__33579));
    LocalMux I__6654 (
            .O(N__33579),
            .I(\delay_measurement_inst.delay_tr_timer.N_320_4 ));
    CascadeMux I__6653 (
            .O(N__33576),
            .I(\delay_measurement_inst.N_305_1_cascade_ ));
    CascadeMux I__6652 (
            .O(N__33573),
            .I(N__33568));
    InMux I__6651 (
            .O(N__33572),
            .I(N__33558));
    InMux I__6650 (
            .O(N__33571),
            .I(N__33558));
    InMux I__6649 (
            .O(N__33568),
            .I(N__33558));
    InMux I__6648 (
            .O(N__33567),
            .I(N__33558));
    LocalMux I__6647 (
            .O(N__33558),
            .I(\delay_measurement_inst.N_305_1 ));
    InMux I__6646 (
            .O(N__33555),
            .I(N__33551));
    InMux I__6645 (
            .O(N__33554),
            .I(N__33548));
    LocalMux I__6644 (
            .O(N__33551),
            .I(N__33545));
    LocalMux I__6643 (
            .O(N__33548),
            .I(\delay_measurement_inst.delay_tr_timer.N_299 ));
    Odrv12 I__6642 (
            .O(N__33545),
            .I(\delay_measurement_inst.delay_tr_timer.N_299 ));
    CascadeMux I__6641 (
            .O(N__33540),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5_cascade_ ));
    CascadeMux I__6640 (
            .O(N__33537),
            .I(\delay_measurement_inst.delay_tr_timer.N_321_cascade_ ));
    CascadeMux I__6639 (
            .O(N__33534),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_ ));
    InMux I__6638 (
            .O(N__33531),
            .I(N__33528));
    LocalMux I__6637 (
            .O(N__33528),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7 ));
    InMux I__6636 (
            .O(N__33525),
            .I(N__33522));
    LocalMux I__6635 (
            .O(N__33522),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ));
    CascadeMux I__6634 (
            .O(N__33519),
            .I(N__33516));
    InMux I__6633 (
            .O(N__33516),
            .I(N__33513));
    LocalMux I__6632 (
            .O(N__33513),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3 ));
    InMux I__6631 (
            .O(N__33510),
            .I(N__33507));
    LocalMux I__6630 (
            .O(N__33507),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ));
    InMux I__6629 (
            .O(N__33504),
            .I(N__33501));
    LocalMux I__6628 (
            .O(N__33501),
            .I(N__33498));
    Span4Mux_h I__6627 (
            .O(N__33498),
            .I(N__33495));
    Odrv4 I__6626 (
            .O(N__33495),
            .I(\current_shift_inst.un4_control_input_axb_12 ));
    InMux I__6625 (
            .O(N__33492),
            .I(N__33489));
    LocalMux I__6624 (
            .O(N__33489),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ));
    InMux I__6623 (
            .O(N__33486),
            .I(N__33483));
    LocalMux I__6622 (
            .O(N__33483),
            .I(N__33480));
    Span4Mux_h I__6621 (
            .O(N__33480),
            .I(N__33477));
    Odrv4 I__6620 (
            .O(N__33477),
            .I(\current_shift_inst.un4_control_input_axb_18 ));
    InMux I__6619 (
            .O(N__33474),
            .I(N__33471));
    LocalMux I__6618 (
            .O(N__33471),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ));
    InMux I__6617 (
            .O(N__33468),
            .I(N__33465));
    LocalMux I__6616 (
            .O(N__33465),
            .I(N__33462));
    Span4Mux_v I__6615 (
            .O(N__33462),
            .I(N__33459));
    Odrv4 I__6614 (
            .O(N__33459),
            .I(\current_shift_inst.un4_control_input_axb_13 ));
    InMux I__6613 (
            .O(N__33456),
            .I(N__33453));
    LocalMux I__6612 (
            .O(N__33453),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ));
    InMux I__6611 (
            .O(N__33450),
            .I(N__33447));
    LocalMux I__6610 (
            .O(N__33447),
            .I(N__33444));
    Span4Mux_h I__6609 (
            .O(N__33444),
            .I(N__33441));
    Odrv4 I__6608 (
            .O(N__33441),
            .I(\current_shift_inst.un4_control_input_axb_14 ));
    InMux I__6607 (
            .O(N__33438),
            .I(N__33435));
    LocalMux I__6606 (
            .O(N__33435),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ));
    InMux I__6605 (
            .O(N__33432),
            .I(N__33429));
    LocalMux I__6604 (
            .O(N__33429),
            .I(N__33426));
    Span4Mux_h I__6603 (
            .O(N__33426),
            .I(N__33423));
    Odrv4 I__6602 (
            .O(N__33423),
            .I(\current_shift_inst.un4_control_input_axb_23 ));
    InMux I__6601 (
            .O(N__33420),
            .I(N__33417));
    LocalMux I__6600 (
            .O(N__33417),
            .I(N__33414));
    Span4Mux_v I__6599 (
            .O(N__33414),
            .I(N__33411));
    Odrv4 I__6598 (
            .O(N__33411),
            .I(\current_shift_inst.un4_control_input_axb_15 ));
    InMux I__6597 (
            .O(N__33408),
            .I(N__33405));
    LocalMux I__6596 (
            .O(N__33405),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ));
    InMux I__6595 (
            .O(N__33402),
            .I(N__33399));
    LocalMux I__6594 (
            .O(N__33399),
            .I(N__33396));
    Span4Mux_h I__6593 (
            .O(N__33396),
            .I(N__33393));
    Odrv4 I__6592 (
            .O(N__33393),
            .I(\current_shift_inst.un4_control_input_axb_16 ));
    InMux I__6591 (
            .O(N__33390),
            .I(N__33387));
    LocalMux I__6590 (
            .O(N__33387),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ));
    InMux I__6589 (
            .O(N__33384),
            .I(N__33381));
    LocalMux I__6588 (
            .O(N__33381),
            .I(N__33378));
    Span4Mux_v I__6587 (
            .O(N__33378),
            .I(N__33375));
    Odrv4 I__6586 (
            .O(N__33375),
            .I(\current_shift_inst.un4_control_input_axb_17 ));
    InMux I__6585 (
            .O(N__33372),
            .I(N__33366));
    InMux I__6584 (
            .O(N__33371),
            .I(N__33361));
    InMux I__6583 (
            .O(N__33370),
            .I(N__33361));
    InMux I__6582 (
            .O(N__33369),
            .I(N__33358));
    LocalMux I__6581 (
            .O(N__33366),
            .I(N__33355));
    LocalMux I__6580 (
            .O(N__33361),
            .I(N__33352));
    LocalMux I__6579 (
            .O(N__33358),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__6578 (
            .O(N__33355),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__6577 (
            .O(N__33352),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__6576 (
            .O(N__33345),
            .I(N__33323));
    InMux I__6575 (
            .O(N__33344),
            .I(N__33323));
    InMux I__6574 (
            .O(N__33343),
            .I(N__33323));
    InMux I__6573 (
            .O(N__33342),
            .I(N__33323));
    InMux I__6572 (
            .O(N__33341),
            .I(N__33302));
    InMux I__6571 (
            .O(N__33340),
            .I(N__33302));
    InMux I__6570 (
            .O(N__33339),
            .I(N__33293));
    InMux I__6569 (
            .O(N__33338),
            .I(N__33293));
    InMux I__6568 (
            .O(N__33337),
            .I(N__33293));
    InMux I__6567 (
            .O(N__33336),
            .I(N__33293));
    InMux I__6566 (
            .O(N__33335),
            .I(N__33284));
    InMux I__6565 (
            .O(N__33334),
            .I(N__33284));
    InMux I__6564 (
            .O(N__33333),
            .I(N__33284));
    InMux I__6563 (
            .O(N__33332),
            .I(N__33284));
    LocalMux I__6562 (
            .O(N__33323),
            .I(N__33281));
    InMux I__6561 (
            .O(N__33322),
            .I(N__33272));
    InMux I__6560 (
            .O(N__33321),
            .I(N__33272));
    InMux I__6559 (
            .O(N__33320),
            .I(N__33272));
    InMux I__6558 (
            .O(N__33319),
            .I(N__33272));
    InMux I__6557 (
            .O(N__33318),
            .I(N__33263));
    InMux I__6556 (
            .O(N__33317),
            .I(N__33263));
    InMux I__6555 (
            .O(N__33316),
            .I(N__33263));
    InMux I__6554 (
            .O(N__33315),
            .I(N__33263));
    InMux I__6553 (
            .O(N__33314),
            .I(N__33254));
    InMux I__6552 (
            .O(N__33313),
            .I(N__33254));
    InMux I__6551 (
            .O(N__33312),
            .I(N__33254));
    InMux I__6550 (
            .O(N__33311),
            .I(N__33254));
    InMux I__6549 (
            .O(N__33310),
            .I(N__33245));
    InMux I__6548 (
            .O(N__33309),
            .I(N__33245));
    InMux I__6547 (
            .O(N__33308),
            .I(N__33245));
    InMux I__6546 (
            .O(N__33307),
            .I(N__33245));
    LocalMux I__6545 (
            .O(N__33302),
            .I(N__33242));
    LocalMux I__6544 (
            .O(N__33293),
            .I(N__33239));
    LocalMux I__6543 (
            .O(N__33284),
            .I(N__33236));
    Span4Mux_h I__6542 (
            .O(N__33281),
            .I(N__33221));
    LocalMux I__6541 (
            .O(N__33272),
            .I(N__33221));
    LocalMux I__6540 (
            .O(N__33263),
            .I(N__33221));
    LocalMux I__6539 (
            .O(N__33254),
            .I(N__33221));
    LocalMux I__6538 (
            .O(N__33245),
            .I(N__33221));
    Span4Mux_v I__6537 (
            .O(N__33242),
            .I(N__33221));
    Span4Mux_v I__6536 (
            .O(N__33239),
            .I(N__33221));
    Span4Mux_v I__6535 (
            .O(N__33236),
            .I(N__33216));
    Span4Mux_v I__6534 (
            .O(N__33221),
            .I(N__33216));
    Odrv4 I__6533 (
            .O(N__33216),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__6532 (
            .O(N__33213),
            .I(N__33210));
    LocalMux I__6531 (
            .O(N__33210),
            .I(N__33207));
    Odrv4 I__6530 (
            .O(N__33207),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ));
    InMux I__6529 (
            .O(N__33204),
            .I(N__33201));
    LocalMux I__6528 (
            .O(N__33201),
            .I(N__33198));
    Span4Mux_v I__6527 (
            .O(N__33198),
            .I(N__33195));
    Odrv4 I__6526 (
            .O(N__33195),
            .I(\current_shift_inst.un4_control_input_axb_21 ));
    InMux I__6525 (
            .O(N__33192),
            .I(N__33189));
    LocalMux I__6524 (
            .O(N__33189),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ));
    InMux I__6523 (
            .O(N__33186),
            .I(N__33183));
    LocalMux I__6522 (
            .O(N__33183),
            .I(N__33180));
    Span4Mux_v I__6521 (
            .O(N__33180),
            .I(N__33177));
    Odrv4 I__6520 (
            .O(N__33177),
            .I(\current_shift_inst.un4_control_input_axb_10 ));
    InMux I__6519 (
            .O(N__33174),
            .I(N__33171));
    LocalMux I__6518 (
            .O(N__33171),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ));
    InMux I__6517 (
            .O(N__33168),
            .I(N__33165));
    LocalMux I__6516 (
            .O(N__33165),
            .I(N__33162));
    Span4Mux_v I__6515 (
            .O(N__33162),
            .I(N__33159));
    Odrv4 I__6514 (
            .O(N__33159),
            .I(\current_shift_inst.un4_control_input_axb_11 ));
    CascadeMux I__6513 (
            .O(N__33156),
            .I(N__33151));
    CascadeMux I__6512 (
            .O(N__33155),
            .I(N__33148));
    InMux I__6511 (
            .O(N__33154),
            .I(N__33145));
    InMux I__6510 (
            .O(N__33151),
            .I(N__33142));
    InMux I__6509 (
            .O(N__33148),
            .I(N__33137));
    LocalMux I__6508 (
            .O(N__33145),
            .I(N__33134));
    LocalMux I__6507 (
            .O(N__33142),
            .I(N__33131));
    InMux I__6506 (
            .O(N__33141),
            .I(N__33126));
    InMux I__6505 (
            .O(N__33140),
            .I(N__33126));
    LocalMux I__6504 (
            .O(N__33137),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__6503 (
            .O(N__33134),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__6502 (
            .O(N__33131),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__6501 (
            .O(N__33126),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__6500 (
            .O(N__33117),
            .I(N__33111));
    InMux I__6499 (
            .O(N__33116),
            .I(N__33108));
    InMux I__6498 (
            .O(N__33115),
            .I(N__33103));
    InMux I__6497 (
            .O(N__33114),
            .I(N__33103));
    LocalMux I__6496 (
            .O(N__33111),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6495 (
            .O(N__33108),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6494 (
            .O(N__33103),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    InMux I__6493 (
            .O(N__33096),
            .I(N__33092));
    InMux I__6492 (
            .O(N__33095),
            .I(N__33089));
    LocalMux I__6491 (
            .O(N__33092),
            .I(N__33085));
    LocalMux I__6490 (
            .O(N__33089),
            .I(N__33082));
    InMux I__6489 (
            .O(N__33088),
            .I(N__33079));
    Odrv4 I__6488 (
            .O(N__33085),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    Odrv4 I__6487 (
            .O(N__33082),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__6486 (
            .O(N__33079),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    InMux I__6485 (
            .O(N__33072),
            .I(N__33069));
    LocalMux I__6484 (
            .O(N__33069),
            .I(N__33065));
    InMux I__6483 (
            .O(N__33068),
            .I(N__33062));
    Span4Mux_h I__6482 (
            .O(N__33065),
            .I(N__33058));
    LocalMux I__6481 (
            .O(N__33062),
            .I(N__33055));
    InMux I__6480 (
            .O(N__33061),
            .I(N__33052));
    Odrv4 I__6479 (
            .O(N__33058),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    Odrv4 I__6478 (
            .O(N__33055),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__6477 (
            .O(N__33052),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    InMux I__6476 (
            .O(N__33045),
            .I(N__33041));
    InMux I__6475 (
            .O(N__33044),
            .I(N__33037));
    LocalMux I__6474 (
            .O(N__33041),
            .I(N__33034));
    InMux I__6473 (
            .O(N__33040),
            .I(N__33031));
    LocalMux I__6472 (
            .O(N__33037),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    Odrv4 I__6471 (
            .O(N__33034),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__6470 (
            .O(N__33031),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    CEMux I__6469 (
            .O(N__33024),
            .I(N__33021));
    LocalMux I__6468 (
            .O(N__33021),
            .I(N__33018));
    Sp12to4 I__6467 (
            .O(N__33018),
            .I(N__33015));
    Odrv12 I__6466 (
            .O(N__33015),
            .I(\phase_controller_inst1.N_221_0 ));
    InMux I__6465 (
            .O(N__33012),
            .I(N__33006));
    InMux I__6464 (
            .O(N__33011),
            .I(N__33006));
    LocalMux I__6463 (
            .O(N__33006),
            .I(N__33003));
    Odrv4 I__6462 (
            .O(N__33003),
            .I(\current_shift_inst.S3_syncZ0Z1 ));
    InMux I__6461 (
            .O(N__33000),
            .I(N__32997));
    LocalMux I__6460 (
            .O(N__32997),
            .I(\current_shift_inst.S3_syncZ0Z0 ));
    InMux I__6459 (
            .O(N__32994),
            .I(N__32991));
    LocalMux I__6458 (
            .O(N__32991),
            .I(N__32988));
    Odrv4 I__6457 (
            .O(N__32988),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ));
    InMux I__6456 (
            .O(N__32985),
            .I(N__32982));
    LocalMux I__6455 (
            .O(N__32982),
            .I(N__32979));
    Span4Mux_v I__6454 (
            .O(N__32979),
            .I(N__32976));
    Odrv4 I__6453 (
            .O(N__32976),
            .I(\current_shift_inst.un4_control_input_axb_24 ));
    InMux I__6452 (
            .O(N__32973),
            .I(N__32970));
    LocalMux I__6451 (
            .O(N__32970),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ));
    CascadeMux I__6450 (
            .O(N__32967),
            .I(N__32963));
    InMux I__6449 (
            .O(N__32966),
            .I(N__32960));
    InMux I__6448 (
            .O(N__32963),
            .I(N__32957));
    LocalMux I__6447 (
            .O(N__32960),
            .I(N__32954));
    LocalMux I__6446 (
            .O(N__32957),
            .I(measured_delay_hc_26));
    Odrv4 I__6445 (
            .O(N__32954),
            .I(measured_delay_hc_26));
    InMux I__6444 (
            .O(N__32949),
            .I(N__32945));
    InMux I__6443 (
            .O(N__32948),
            .I(N__32942));
    LocalMux I__6442 (
            .O(N__32945),
            .I(N__32939));
    LocalMux I__6441 (
            .O(N__32942),
            .I(measured_delay_hc_24));
    Odrv4 I__6440 (
            .O(N__32939),
            .I(measured_delay_hc_24));
    IoInMux I__6439 (
            .O(N__32934),
            .I(N__32931));
    LocalMux I__6438 (
            .O(N__32931),
            .I(N__32928));
    IoSpan4Mux I__6437 (
            .O(N__32928),
            .I(N__32925));
    Span4Mux_s1_v I__6436 (
            .O(N__32925),
            .I(N__32921));
    InMux I__6435 (
            .O(N__32924),
            .I(N__32918));
    Sp12to4 I__6434 (
            .O(N__32921),
            .I(N__32915));
    LocalMux I__6433 (
            .O(N__32918),
            .I(N__32912));
    Span12Mux_s8_v I__6432 (
            .O(N__32915),
            .I(N__32909));
    Span4Mux_v I__6431 (
            .O(N__32912),
            .I(N__32906));
    Odrv12 I__6430 (
            .O(N__32909),
            .I(s1_phy_c));
    Odrv4 I__6429 (
            .O(N__32906),
            .I(s1_phy_c));
    InMux I__6428 (
            .O(N__32901),
            .I(N__32898));
    LocalMux I__6427 (
            .O(N__32898),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ));
    InMux I__6426 (
            .O(N__32895),
            .I(N__32891));
    CascadeMux I__6425 (
            .O(N__32894),
            .I(N__32888));
    LocalMux I__6424 (
            .O(N__32891),
            .I(N__32885));
    InMux I__6423 (
            .O(N__32888),
            .I(N__32882));
    Span4Mux_h I__6422 (
            .O(N__32885),
            .I(N__32879));
    LocalMux I__6421 (
            .O(N__32882),
            .I(measured_delay_hc_25));
    Odrv4 I__6420 (
            .O(N__32879),
            .I(measured_delay_hc_25));
    InMux I__6419 (
            .O(N__32874),
            .I(N__32840));
    InMux I__6418 (
            .O(N__32873),
            .I(N__32840));
    InMux I__6417 (
            .O(N__32872),
            .I(N__32840));
    InMux I__6416 (
            .O(N__32871),
            .I(N__32840));
    InMux I__6415 (
            .O(N__32870),
            .I(N__32840));
    InMux I__6414 (
            .O(N__32869),
            .I(N__32840));
    InMux I__6413 (
            .O(N__32868),
            .I(N__32840));
    InMux I__6412 (
            .O(N__32867),
            .I(N__32825));
    InMux I__6411 (
            .O(N__32866),
            .I(N__32825));
    InMux I__6410 (
            .O(N__32865),
            .I(N__32825));
    InMux I__6409 (
            .O(N__32864),
            .I(N__32825));
    InMux I__6408 (
            .O(N__32863),
            .I(N__32825));
    InMux I__6407 (
            .O(N__32862),
            .I(N__32825));
    InMux I__6406 (
            .O(N__32861),
            .I(N__32825));
    InMux I__6405 (
            .O(N__32860),
            .I(N__32814));
    InMux I__6404 (
            .O(N__32859),
            .I(N__32814));
    InMux I__6403 (
            .O(N__32858),
            .I(N__32814));
    InMux I__6402 (
            .O(N__32857),
            .I(N__32814));
    InMux I__6401 (
            .O(N__32856),
            .I(N__32814));
    InMux I__6400 (
            .O(N__32855),
            .I(N__32809));
    LocalMux I__6399 (
            .O(N__32840),
            .I(N__32804));
    LocalMux I__6398 (
            .O(N__32825),
            .I(N__32804));
    LocalMux I__6397 (
            .O(N__32814),
            .I(N__32800));
    InMux I__6396 (
            .O(N__32813),
            .I(N__32797));
    InMux I__6395 (
            .O(N__32812),
            .I(N__32793));
    LocalMux I__6394 (
            .O(N__32809),
            .I(N__32790));
    Span4Mux_v I__6393 (
            .O(N__32804),
            .I(N__32787));
    InMux I__6392 (
            .O(N__32803),
            .I(N__32784));
    Span4Mux_h I__6391 (
            .O(N__32800),
            .I(N__32779));
    LocalMux I__6390 (
            .O(N__32797),
            .I(N__32779));
    InMux I__6389 (
            .O(N__32796),
            .I(N__32776));
    LocalMux I__6388 (
            .O(N__32793),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__6387 (
            .O(N__32790),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__6386 (
            .O(N__32787),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__6385 (
            .O(N__32784),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__6384 (
            .O(N__32779),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__6383 (
            .O(N__32776),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__6382 (
            .O(N__32763),
            .I(N__32757));
    CascadeMux I__6381 (
            .O(N__32762),
            .I(N__32754));
    CascadeMux I__6380 (
            .O(N__32761),
            .I(N__32751));
    InMux I__6379 (
            .O(N__32760),
            .I(N__32732));
    InMux I__6378 (
            .O(N__32757),
            .I(N__32722));
    InMux I__6377 (
            .O(N__32754),
            .I(N__32722));
    InMux I__6376 (
            .O(N__32751),
            .I(N__32722));
    InMux I__6375 (
            .O(N__32750),
            .I(N__32719));
    InMux I__6374 (
            .O(N__32749),
            .I(N__32704));
    InMux I__6373 (
            .O(N__32748),
            .I(N__32704));
    InMux I__6372 (
            .O(N__32747),
            .I(N__32704));
    InMux I__6371 (
            .O(N__32746),
            .I(N__32704));
    InMux I__6370 (
            .O(N__32745),
            .I(N__32704));
    InMux I__6369 (
            .O(N__32744),
            .I(N__32704));
    InMux I__6368 (
            .O(N__32743),
            .I(N__32704));
    InMux I__6367 (
            .O(N__32742),
            .I(N__32689));
    InMux I__6366 (
            .O(N__32741),
            .I(N__32689));
    InMux I__6365 (
            .O(N__32740),
            .I(N__32689));
    InMux I__6364 (
            .O(N__32739),
            .I(N__32689));
    InMux I__6363 (
            .O(N__32738),
            .I(N__32689));
    InMux I__6362 (
            .O(N__32737),
            .I(N__32689));
    InMux I__6361 (
            .O(N__32736),
            .I(N__32689));
    InMux I__6360 (
            .O(N__32735),
            .I(N__32686));
    LocalMux I__6359 (
            .O(N__32732),
            .I(N__32683));
    InMux I__6358 (
            .O(N__32731),
            .I(N__32679));
    InMux I__6357 (
            .O(N__32730),
            .I(N__32674));
    InMux I__6356 (
            .O(N__32729),
            .I(N__32674));
    LocalMux I__6355 (
            .O(N__32722),
            .I(N__32669));
    LocalMux I__6354 (
            .O(N__32719),
            .I(N__32669));
    LocalMux I__6353 (
            .O(N__32704),
            .I(N__32666));
    LocalMux I__6352 (
            .O(N__32689),
            .I(N__32663));
    LocalMux I__6351 (
            .O(N__32686),
            .I(N__32658));
    Span4Mux_v I__6350 (
            .O(N__32683),
            .I(N__32658));
    InMux I__6349 (
            .O(N__32682),
            .I(N__32655));
    LocalMux I__6348 (
            .O(N__32679),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__6347 (
            .O(N__32674),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__6346 (
            .O(N__32669),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__6345 (
            .O(N__32666),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__6344 (
            .O(N__32663),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__6343 (
            .O(N__32658),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__6342 (
            .O(N__32655),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    InMux I__6341 (
            .O(N__32640),
            .I(N__32637));
    LocalMux I__6340 (
            .O(N__32637),
            .I(N__32634));
    Glb2LocalMux I__6339 (
            .O(N__32634),
            .I(N__32631));
    GlobalMux I__6338 (
            .O(N__32631),
            .I(clk_12mhz));
    IoInMux I__6337 (
            .O(N__32628),
            .I(N__32625));
    LocalMux I__6336 (
            .O(N__32625),
            .I(N__32622));
    Span4Mux_s0_v I__6335 (
            .O(N__32622),
            .I(N__32619));
    Odrv4 I__6334 (
            .O(N__32619),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__6333 (
            .O(N__32616),
            .I(N__32613));
    LocalMux I__6332 (
            .O(N__32613),
            .I(N__32610));
    Span4Mux_v I__6331 (
            .O(N__32610),
            .I(N__32607));
    Span4Mux_h I__6330 (
            .O(N__32607),
            .I(N__32604));
    Span4Mux_h I__6329 (
            .O(N__32604),
            .I(N__32601));
    Odrv4 I__6328 (
            .O(N__32601),
            .I(il_max_comp2_c));
    InMux I__6327 (
            .O(N__32598),
            .I(N__32595));
    LocalMux I__6326 (
            .O(N__32595),
            .I(il_max_comp2_D1));
    CascadeMux I__6325 (
            .O(N__32592),
            .I(N__32588));
    CascadeMux I__6324 (
            .O(N__32591),
            .I(N__32585));
    InMux I__6323 (
            .O(N__32588),
            .I(N__32580));
    InMux I__6322 (
            .O(N__32585),
            .I(N__32580));
    LocalMux I__6321 (
            .O(N__32580),
            .I(N__32576));
    InMux I__6320 (
            .O(N__32579),
            .I(N__32573));
    Span4Mux_v I__6319 (
            .O(N__32576),
            .I(N__32570));
    LocalMux I__6318 (
            .O(N__32573),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__6317 (
            .O(N__32570),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__6316 (
            .O(N__32565),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__6315 (
            .O(N__32562),
            .I(N__32558));
    InMux I__6314 (
            .O(N__32561),
            .I(N__32555));
    LocalMux I__6313 (
            .O(N__32558),
            .I(N__32549));
    LocalMux I__6312 (
            .O(N__32555),
            .I(N__32549));
    InMux I__6311 (
            .O(N__32554),
            .I(N__32546));
    Span4Mux_v I__6310 (
            .O(N__32549),
            .I(N__32543));
    LocalMux I__6309 (
            .O(N__32546),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__6308 (
            .O(N__32543),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__6307 (
            .O(N__32538),
            .I(bfn_12_22_0_));
    CascadeMux I__6306 (
            .O(N__32535),
            .I(N__32532));
    InMux I__6305 (
            .O(N__32532),
            .I(N__32528));
    InMux I__6304 (
            .O(N__32531),
            .I(N__32525));
    LocalMux I__6303 (
            .O(N__32528),
            .I(N__32519));
    LocalMux I__6302 (
            .O(N__32525),
            .I(N__32519));
    InMux I__6301 (
            .O(N__32524),
            .I(N__32516));
    Span4Mux_v I__6300 (
            .O(N__32519),
            .I(N__32513));
    LocalMux I__6299 (
            .O(N__32516),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__6298 (
            .O(N__32513),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__6297 (
            .O(N__32508),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__6296 (
            .O(N__32505),
            .I(N__32501));
    CascadeMux I__6295 (
            .O(N__32504),
            .I(N__32498));
    InMux I__6294 (
            .O(N__32501),
            .I(N__32493));
    InMux I__6293 (
            .O(N__32498),
            .I(N__32493));
    LocalMux I__6292 (
            .O(N__32493),
            .I(N__32489));
    InMux I__6291 (
            .O(N__32492),
            .I(N__32486));
    Span4Mux_v I__6290 (
            .O(N__32489),
            .I(N__32483));
    LocalMux I__6289 (
            .O(N__32486),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__6288 (
            .O(N__32483),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__6287 (
            .O(N__32478),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__6286 (
            .O(N__32475),
            .I(N__32468));
    InMux I__6285 (
            .O(N__32474),
            .I(N__32468));
    InMux I__6284 (
            .O(N__32473),
            .I(N__32465));
    LocalMux I__6283 (
            .O(N__32468),
            .I(N__32462));
    LocalMux I__6282 (
            .O(N__32465),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv12 I__6281 (
            .O(N__32462),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__6280 (
            .O(N__32457),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__6279 (
            .O(N__32454),
            .I(N__32451));
    LocalMux I__6278 (
            .O(N__32451),
            .I(N__32447));
    InMux I__6277 (
            .O(N__32450),
            .I(N__32444));
    Span4Mux_v I__6276 (
            .O(N__32447),
            .I(N__32441));
    LocalMux I__6275 (
            .O(N__32444),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__6274 (
            .O(N__32441),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__6273 (
            .O(N__32436),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__6272 (
            .O(N__32433),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CascadeMux I__6271 (
            .O(N__32430),
            .I(N__32427));
    InMux I__6270 (
            .O(N__32427),
            .I(N__32423));
    InMux I__6269 (
            .O(N__32426),
            .I(N__32420));
    LocalMux I__6268 (
            .O(N__32423),
            .I(N__32417));
    LocalMux I__6267 (
            .O(N__32420),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv12 I__6266 (
            .O(N__32417),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__6265 (
            .O(N__32412),
            .I(N__32408));
    CEMux I__6264 (
            .O(N__32411),
            .I(N__32405));
    LocalMux I__6263 (
            .O(N__32408),
            .I(N__32398));
    LocalMux I__6262 (
            .O(N__32405),
            .I(N__32398));
    CEMux I__6261 (
            .O(N__32404),
            .I(N__32395));
    CEMux I__6260 (
            .O(N__32403),
            .I(N__32392));
    Span4Mux_v I__6259 (
            .O(N__32398),
            .I(N__32389));
    LocalMux I__6258 (
            .O(N__32395),
            .I(N__32384));
    LocalMux I__6257 (
            .O(N__32392),
            .I(N__32384));
    Span4Mux_h I__6256 (
            .O(N__32389),
            .I(N__32379));
    Span4Mux_v I__6255 (
            .O(N__32384),
            .I(N__32379));
    Span4Mux_v I__6254 (
            .O(N__32379),
            .I(N__32376));
    Odrv4 I__6253 (
            .O(N__32376),
            .I(\current_shift_inst.timer_s1.N_191_i ));
    IoInMux I__6252 (
            .O(N__32373),
            .I(N__32370));
    LocalMux I__6251 (
            .O(N__32370),
            .I(N__32367));
    Span4Mux_s0_v I__6250 (
            .O(N__32367),
            .I(N__32364));
    Span4Mux_v I__6249 (
            .O(N__32364),
            .I(N__32361));
    Odrv4 I__6248 (
            .O(N__32361),
            .I(\current_shift_inst.timer_phase.N_188_i ));
    CascadeMux I__6247 (
            .O(N__32358),
            .I(N__32354));
    CascadeMux I__6246 (
            .O(N__32357),
            .I(N__32351));
    InMux I__6245 (
            .O(N__32354),
            .I(N__32346));
    InMux I__6244 (
            .O(N__32351),
            .I(N__32346));
    LocalMux I__6243 (
            .O(N__32346),
            .I(N__32342));
    InMux I__6242 (
            .O(N__32345),
            .I(N__32339));
    Span4Mux_v I__6241 (
            .O(N__32342),
            .I(N__32336));
    LocalMux I__6240 (
            .O(N__32339),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__6239 (
            .O(N__32336),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__6238 (
            .O(N__32331),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__6237 (
            .O(N__32328),
            .I(N__32324));
    InMux I__6236 (
            .O(N__32327),
            .I(N__32321));
    InMux I__6235 (
            .O(N__32324),
            .I(N__32318));
    LocalMux I__6234 (
            .O(N__32321),
            .I(N__32312));
    LocalMux I__6233 (
            .O(N__32318),
            .I(N__32312));
    InMux I__6232 (
            .O(N__32317),
            .I(N__32309));
    Span4Mux_v I__6231 (
            .O(N__32312),
            .I(N__32306));
    LocalMux I__6230 (
            .O(N__32309),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__6229 (
            .O(N__32306),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__6228 (
            .O(N__32301),
            .I(bfn_12_21_0_));
    InMux I__6227 (
            .O(N__32298),
            .I(N__32294));
    InMux I__6226 (
            .O(N__32297),
            .I(N__32291));
    LocalMux I__6225 (
            .O(N__32294),
            .I(N__32285));
    LocalMux I__6224 (
            .O(N__32291),
            .I(N__32285));
    InMux I__6223 (
            .O(N__32290),
            .I(N__32282));
    Span4Mux_v I__6222 (
            .O(N__32285),
            .I(N__32279));
    LocalMux I__6221 (
            .O(N__32282),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__6220 (
            .O(N__32279),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__6219 (
            .O(N__32274),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    CascadeMux I__6218 (
            .O(N__32271),
            .I(N__32267));
    CascadeMux I__6217 (
            .O(N__32270),
            .I(N__32264));
    InMux I__6216 (
            .O(N__32267),
            .I(N__32259));
    InMux I__6215 (
            .O(N__32264),
            .I(N__32259));
    LocalMux I__6214 (
            .O(N__32259),
            .I(N__32255));
    InMux I__6213 (
            .O(N__32258),
            .I(N__32252));
    Span4Mux_v I__6212 (
            .O(N__32255),
            .I(N__32249));
    LocalMux I__6211 (
            .O(N__32252),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__6210 (
            .O(N__32249),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__6209 (
            .O(N__32244),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__6208 (
            .O(N__32241),
            .I(N__32237));
    CascadeMux I__6207 (
            .O(N__32240),
            .I(N__32234));
    InMux I__6206 (
            .O(N__32237),
            .I(N__32229));
    InMux I__6205 (
            .O(N__32234),
            .I(N__32229));
    LocalMux I__6204 (
            .O(N__32229),
            .I(N__32225));
    InMux I__6203 (
            .O(N__32228),
            .I(N__32222));
    Span4Mux_v I__6202 (
            .O(N__32225),
            .I(N__32219));
    LocalMux I__6201 (
            .O(N__32222),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__6200 (
            .O(N__32219),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__6199 (
            .O(N__32214),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__6198 (
            .O(N__32211),
            .I(N__32205));
    InMux I__6197 (
            .O(N__32210),
            .I(N__32205));
    LocalMux I__6196 (
            .O(N__32205),
            .I(N__32201));
    InMux I__6195 (
            .O(N__32204),
            .I(N__32198));
    Span4Mux_v I__6194 (
            .O(N__32201),
            .I(N__32195));
    LocalMux I__6193 (
            .O(N__32198),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__6192 (
            .O(N__32195),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__6191 (
            .O(N__32190),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__6190 (
            .O(N__32187),
            .I(N__32180));
    InMux I__6189 (
            .O(N__32186),
            .I(N__32180));
    InMux I__6188 (
            .O(N__32185),
            .I(N__32177));
    LocalMux I__6187 (
            .O(N__32180),
            .I(N__32174));
    LocalMux I__6186 (
            .O(N__32177),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv12 I__6185 (
            .O(N__32174),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__6184 (
            .O(N__32169),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__6183 (
            .O(N__32166),
            .I(N__32162));
    CascadeMux I__6182 (
            .O(N__32165),
            .I(N__32159));
    InMux I__6181 (
            .O(N__32162),
            .I(N__32153));
    InMux I__6180 (
            .O(N__32159),
            .I(N__32153));
    InMux I__6179 (
            .O(N__32158),
            .I(N__32150));
    LocalMux I__6178 (
            .O(N__32153),
            .I(N__32147));
    LocalMux I__6177 (
            .O(N__32150),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv12 I__6176 (
            .O(N__32147),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__6175 (
            .O(N__32142),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__6174 (
            .O(N__32139),
            .I(N__32135));
    CascadeMux I__6173 (
            .O(N__32138),
            .I(N__32132));
    InMux I__6172 (
            .O(N__32135),
            .I(N__32126));
    InMux I__6171 (
            .O(N__32132),
            .I(N__32126));
    InMux I__6170 (
            .O(N__32131),
            .I(N__32123));
    LocalMux I__6169 (
            .O(N__32126),
            .I(N__32120));
    LocalMux I__6168 (
            .O(N__32123),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv12 I__6167 (
            .O(N__32120),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__6166 (
            .O(N__32115),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    CascadeMux I__6165 (
            .O(N__32112),
            .I(N__32108));
    CascadeMux I__6164 (
            .O(N__32111),
            .I(N__32105));
    InMux I__6163 (
            .O(N__32108),
            .I(N__32100));
    InMux I__6162 (
            .O(N__32105),
            .I(N__32100));
    LocalMux I__6161 (
            .O(N__32100),
            .I(N__32096));
    InMux I__6160 (
            .O(N__32099),
            .I(N__32093));
    Span4Mux_v I__6159 (
            .O(N__32096),
            .I(N__32090));
    LocalMux I__6158 (
            .O(N__32093),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__6157 (
            .O(N__32090),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__6156 (
            .O(N__32085),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    InMux I__6155 (
            .O(N__32082),
            .I(N__32078));
    InMux I__6154 (
            .O(N__32081),
            .I(N__32075));
    LocalMux I__6153 (
            .O(N__32078),
            .I(N__32069));
    LocalMux I__6152 (
            .O(N__32075),
            .I(N__32069));
    InMux I__6151 (
            .O(N__32074),
            .I(N__32066));
    Span4Mux_v I__6150 (
            .O(N__32069),
            .I(N__32063));
    LocalMux I__6149 (
            .O(N__32066),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__6148 (
            .O(N__32063),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__6147 (
            .O(N__32058),
            .I(bfn_12_20_0_));
    InMux I__6146 (
            .O(N__32055),
            .I(N__32050));
    InMux I__6145 (
            .O(N__32054),
            .I(N__32047));
    InMux I__6144 (
            .O(N__32053),
            .I(N__32044));
    LocalMux I__6143 (
            .O(N__32050),
            .I(N__32039));
    LocalMux I__6142 (
            .O(N__32047),
            .I(N__32039));
    LocalMux I__6141 (
            .O(N__32044),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv12 I__6140 (
            .O(N__32039),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__6139 (
            .O(N__32034),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__6138 (
            .O(N__32031),
            .I(N__32027));
    CascadeMux I__6137 (
            .O(N__32030),
            .I(N__32024));
    InMux I__6136 (
            .O(N__32027),
            .I(N__32018));
    InMux I__6135 (
            .O(N__32024),
            .I(N__32018));
    InMux I__6134 (
            .O(N__32023),
            .I(N__32015));
    LocalMux I__6133 (
            .O(N__32018),
            .I(N__32012));
    LocalMux I__6132 (
            .O(N__32015),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv12 I__6131 (
            .O(N__32012),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__6130 (
            .O(N__32007),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    CascadeMux I__6129 (
            .O(N__32004),
            .I(N__32000));
    CascadeMux I__6128 (
            .O(N__32003),
            .I(N__31997));
    InMux I__6127 (
            .O(N__32000),
            .I(N__31991));
    InMux I__6126 (
            .O(N__31997),
            .I(N__31991));
    InMux I__6125 (
            .O(N__31996),
            .I(N__31988));
    LocalMux I__6124 (
            .O(N__31991),
            .I(N__31985));
    LocalMux I__6123 (
            .O(N__31988),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv12 I__6122 (
            .O(N__31985),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__6121 (
            .O(N__31980),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__6120 (
            .O(N__31977),
            .I(N__31970));
    InMux I__6119 (
            .O(N__31976),
            .I(N__31970));
    InMux I__6118 (
            .O(N__31975),
            .I(N__31967));
    LocalMux I__6117 (
            .O(N__31970),
            .I(N__31964));
    LocalMux I__6116 (
            .O(N__31967),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv12 I__6115 (
            .O(N__31964),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__6114 (
            .O(N__31959),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    InMux I__6113 (
            .O(N__31956),
            .I(N__31950));
    InMux I__6112 (
            .O(N__31955),
            .I(N__31950));
    LocalMux I__6111 (
            .O(N__31950),
            .I(N__31946));
    InMux I__6110 (
            .O(N__31949),
            .I(N__31943));
    Span4Mux_v I__6109 (
            .O(N__31946),
            .I(N__31940));
    LocalMux I__6108 (
            .O(N__31943),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__6107 (
            .O(N__31940),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__6106 (
            .O(N__31935),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__6105 (
            .O(N__31932),
            .I(N__31929));
    InMux I__6104 (
            .O(N__31929),
            .I(N__31925));
    InMux I__6103 (
            .O(N__31928),
            .I(N__31921));
    LocalMux I__6102 (
            .O(N__31925),
            .I(N__31918));
    InMux I__6101 (
            .O(N__31924),
            .I(N__31915));
    LocalMux I__6100 (
            .O(N__31921),
            .I(N__31912));
    Span4Mux_v I__6099 (
            .O(N__31918),
            .I(N__31909));
    LocalMux I__6098 (
            .O(N__31915),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv12 I__6097 (
            .O(N__31912),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__6096 (
            .O(N__31909),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__6095 (
            .O(N__31902),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__6094 (
            .O(N__31899),
            .I(N__31896));
    LocalMux I__6093 (
            .O(N__31896),
            .I(N__31893));
    Odrv4 I__6092 (
            .O(N__31893),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ));
    InMux I__6091 (
            .O(N__31890),
            .I(N__31887));
    LocalMux I__6090 (
            .O(N__31887),
            .I(\current_shift_inst.un4_control_input_axb_25 ));
    InMux I__6089 (
            .O(N__31884),
            .I(N__31881));
    LocalMux I__6088 (
            .O(N__31881),
            .I(N__31878));
    Odrv4 I__6087 (
            .O(N__31878),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ));
    InMux I__6086 (
            .O(N__31875),
            .I(N__31872));
    LocalMux I__6085 (
            .O(N__31872),
            .I(\current_shift_inst.un4_control_input_axb_22 ));
    InMux I__6084 (
            .O(N__31869),
            .I(N__31865));
    CascadeMux I__6083 (
            .O(N__31868),
            .I(N__31862));
    LocalMux I__6082 (
            .O(N__31865),
            .I(N__31859));
    InMux I__6081 (
            .O(N__31862),
            .I(N__31855));
    Span4Mux_h I__6080 (
            .O(N__31859),
            .I(N__31852));
    InMux I__6079 (
            .O(N__31858),
            .I(N__31849));
    LocalMux I__6078 (
            .O(N__31855),
            .I(N__31846));
    Odrv4 I__6077 (
            .O(N__31852),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__6076 (
            .O(N__31849),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv12 I__6075 (
            .O(N__31846),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__6074 (
            .O(N__31839),
            .I(bfn_12_19_0_));
    InMux I__6073 (
            .O(N__31836),
            .I(N__31832));
    CascadeMux I__6072 (
            .O(N__31835),
            .I(N__31829));
    LocalMux I__6071 (
            .O(N__31832),
            .I(N__31826));
    InMux I__6070 (
            .O(N__31829),
            .I(N__31822));
    Span4Mux_h I__6069 (
            .O(N__31826),
            .I(N__31819));
    InMux I__6068 (
            .O(N__31825),
            .I(N__31816));
    LocalMux I__6067 (
            .O(N__31822),
            .I(N__31813));
    Odrv4 I__6066 (
            .O(N__31819),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__6065 (
            .O(N__31816),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv12 I__6064 (
            .O(N__31813),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__6063 (
            .O(N__31806),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__6062 (
            .O(N__31803),
            .I(N__31796));
    InMux I__6061 (
            .O(N__31802),
            .I(N__31796));
    InMux I__6060 (
            .O(N__31801),
            .I(N__31793));
    LocalMux I__6059 (
            .O(N__31796),
            .I(N__31790));
    LocalMux I__6058 (
            .O(N__31793),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__6057 (
            .O(N__31790),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__6056 (
            .O(N__31785),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__6055 (
            .O(N__31782),
            .I(N__31775));
    InMux I__6054 (
            .O(N__31781),
            .I(N__31775));
    InMux I__6053 (
            .O(N__31780),
            .I(N__31772));
    LocalMux I__6052 (
            .O(N__31775),
            .I(N__31769));
    LocalMux I__6051 (
            .O(N__31772),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv12 I__6050 (
            .O(N__31769),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__6049 (
            .O(N__31764),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__6048 (
            .O(N__31761),
            .I(N__31758));
    InMux I__6047 (
            .O(N__31758),
            .I(N__31754));
    InMux I__6046 (
            .O(N__31757),
            .I(N__31750));
    LocalMux I__6045 (
            .O(N__31754),
            .I(N__31747));
    InMux I__6044 (
            .O(N__31753),
            .I(N__31744));
    LocalMux I__6043 (
            .O(N__31750),
            .I(N__31739));
    Sp12to4 I__6042 (
            .O(N__31747),
            .I(N__31739));
    LocalMux I__6041 (
            .O(N__31744),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv12 I__6040 (
            .O(N__31739),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__6039 (
            .O(N__31734),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__6038 (
            .O(N__31731),
            .I(N__31728));
    InMux I__6037 (
            .O(N__31728),
            .I(N__31724));
    InMux I__6036 (
            .O(N__31727),
            .I(N__31720));
    LocalMux I__6035 (
            .O(N__31724),
            .I(N__31717));
    InMux I__6034 (
            .O(N__31723),
            .I(N__31714));
    LocalMux I__6033 (
            .O(N__31720),
            .I(N__31709));
    Sp12to4 I__6032 (
            .O(N__31717),
            .I(N__31709));
    LocalMux I__6031 (
            .O(N__31714),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv12 I__6030 (
            .O(N__31709),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__6029 (
            .O(N__31704),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__6028 (
            .O(N__31701),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    CEMux I__6027 (
            .O(N__31698),
            .I(N__31683));
    CEMux I__6026 (
            .O(N__31697),
            .I(N__31683));
    CEMux I__6025 (
            .O(N__31696),
            .I(N__31683));
    CEMux I__6024 (
            .O(N__31695),
            .I(N__31683));
    CEMux I__6023 (
            .O(N__31694),
            .I(N__31683));
    GlobalMux I__6022 (
            .O(N__31683),
            .I(N__31680));
    gio2CtrlBuf I__6021 (
            .O(N__31680),
            .I(\current_shift_inst.timer_s1.N_187_i_g ));
    InMux I__6020 (
            .O(N__31677),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__6019 (
            .O(N__31674),
            .I(N__31668));
    InMux I__6018 (
            .O(N__31673),
            .I(N__31668));
    LocalMux I__6017 (
            .O(N__31668),
            .I(N__31665));
    Span4Mux_h I__6016 (
            .O(N__31665),
            .I(N__31662));
    Odrv4 I__6015 (
            .O(N__31662),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__6014 (
            .O(N__31659),
            .I(N__31656));
    LocalMux I__6013 (
            .O(N__31656),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ));
    InMux I__6012 (
            .O(N__31653),
            .I(N__31650));
    LocalMux I__6011 (
            .O(N__31650),
            .I(N__31647));
    Odrv4 I__6010 (
            .O(N__31647),
            .I(\current_shift_inst.un4_control_input_axb_29 ));
    InMux I__6009 (
            .O(N__31644),
            .I(N__31641));
    LocalMux I__6008 (
            .O(N__31641),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ));
    InMux I__6007 (
            .O(N__31638),
            .I(N__31635));
    LocalMux I__6006 (
            .O(N__31635),
            .I(\current_shift_inst.un4_control_input_axb_28 ));
    InMux I__6005 (
            .O(N__31632),
            .I(N__31629));
    LocalMux I__6004 (
            .O(N__31629),
            .I(N__31626));
    Odrv4 I__6003 (
            .O(N__31626),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ));
    InMux I__6002 (
            .O(N__31623),
            .I(N__31620));
    LocalMux I__6001 (
            .O(N__31620),
            .I(\current_shift_inst.un4_control_input_axb_20 ));
    InMux I__6000 (
            .O(N__31617),
            .I(N__31614));
    LocalMux I__5999 (
            .O(N__31614),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ));
    CascadeMux I__5998 (
            .O(N__31611),
            .I(N__31608));
    InMux I__5997 (
            .O(N__31608),
            .I(N__31605));
    LocalMux I__5996 (
            .O(N__31605),
            .I(\current_shift_inst.un4_control_input_axb_30 ));
    InMux I__5995 (
            .O(N__31602),
            .I(N__31599));
    LocalMux I__5994 (
            .O(N__31599),
            .I(N__31596));
    Odrv4 I__5993 (
            .O(N__31596),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ));
    CascadeMux I__5992 (
            .O(N__31593),
            .I(N__31590));
    InMux I__5991 (
            .O(N__31590),
            .I(N__31587));
    LocalMux I__5990 (
            .O(N__31587),
            .I(\current_shift_inst.un4_control_input_axb_19 ));
    InMux I__5989 (
            .O(N__31584),
            .I(N__31581));
    LocalMux I__5988 (
            .O(N__31581),
            .I(N__31578));
    Odrv4 I__5987 (
            .O(N__31578),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ));
    InMux I__5986 (
            .O(N__31575),
            .I(N__31572));
    LocalMux I__5985 (
            .O(N__31572),
            .I(\current_shift_inst.un4_control_input_axb_26 ));
    InMux I__5984 (
            .O(N__31569),
            .I(N__31566));
    LocalMux I__5983 (
            .O(N__31566),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ));
    InMux I__5982 (
            .O(N__31563),
            .I(N__31560));
    LocalMux I__5981 (
            .O(N__31560),
            .I(\current_shift_inst.un4_control_input_axb_27 ));
    InMux I__5980 (
            .O(N__31557),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__5979 (
            .O(N__31554),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__5978 (
            .O(N__31551),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__5977 (
            .O(N__31548),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__5976 (
            .O(N__31545),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__5975 (
            .O(N__31542),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__5974 (
            .O(N__31539),
            .I(bfn_12_17_0_));
    InMux I__5973 (
            .O(N__31536),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__5972 (
            .O(N__31533),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__5971 (
            .O(N__31530),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__5970 (
            .O(N__31527),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__5969 (
            .O(N__31524),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__5968 (
            .O(N__31521),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__5967 (
            .O(N__31518),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__5966 (
            .O(N__31515),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__5965 (
            .O(N__31512),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__5964 (
            .O(N__31509),
            .I(bfn_12_16_0_));
    InMux I__5963 (
            .O(N__31506),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__5962 (
            .O(N__31503),
            .I(N__31500));
    LocalMux I__5961 (
            .O(N__31500),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ));
    InMux I__5960 (
            .O(N__31497),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__5959 (
            .O(N__31494),
            .I(N__31491));
    LocalMux I__5958 (
            .O(N__31491),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ));
    InMux I__5957 (
            .O(N__31488),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__5956 (
            .O(N__31485),
            .I(N__31482));
    LocalMux I__5955 (
            .O(N__31482),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ));
    InMux I__5954 (
            .O(N__31479),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__5953 (
            .O(N__31476),
            .I(N__31473));
    LocalMux I__5952 (
            .O(N__31473),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ));
    InMux I__5951 (
            .O(N__31470),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__5950 (
            .O(N__31467),
            .I(N__31464));
    LocalMux I__5949 (
            .O(N__31464),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ));
    InMux I__5948 (
            .O(N__31461),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__5947 (
            .O(N__31458),
            .I(N__31455));
    LocalMux I__5946 (
            .O(N__31455),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ));
    InMux I__5945 (
            .O(N__31452),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__5944 (
            .O(N__31449),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__5943 (
            .O(N__31446),
            .I(bfn_12_15_0_));
    InMux I__5942 (
            .O(N__31443),
            .I(N__31439));
    InMux I__5941 (
            .O(N__31442),
            .I(N__31436));
    LocalMux I__5940 (
            .O(N__31439),
            .I(N__31433));
    LocalMux I__5939 (
            .O(N__31436),
            .I(N__31430));
    Odrv4 I__5938 (
            .O(N__31433),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt15 ));
    Odrv12 I__5937 (
            .O(N__31430),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt15 ));
    InMux I__5936 (
            .O(N__31425),
            .I(N__31422));
    LocalMux I__5935 (
            .O(N__31422),
            .I(N__31417));
    CascadeMux I__5934 (
            .O(N__31421),
            .I(N__31414));
    CascadeMux I__5933 (
            .O(N__31420),
            .I(N__31411));
    Span4Mux_v I__5932 (
            .O(N__31417),
            .I(N__31408));
    InMux I__5931 (
            .O(N__31414),
            .I(N__31405));
    InMux I__5930 (
            .O(N__31411),
            .I(N__31402));
    Odrv4 I__5929 (
            .O(N__31408),
            .I(\current_shift_inst.S3_riseZ0 ));
    LocalMux I__5928 (
            .O(N__31405),
            .I(\current_shift_inst.S3_riseZ0 ));
    LocalMux I__5927 (
            .O(N__31402),
            .I(\current_shift_inst.S3_riseZ0 ));
    InMux I__5926 (
            .O(N__31395),
            .I(N__31389));
    InMux I__5925 (
            .O(N__31394),
            .I(N__31386));
    InMux I__5924 (
            .O(N__31393),
            .I(N__31381));
    InMux I__5923 (
            .O(N__31392),
            .I(N__31381));
    LocalMux I__5922 (
            .O(N__31389),
            .I(N__31374));
    LocalMux I__5921 (
            .O(N__31386),
            .I(N__31374));
    LocalMux I__5920 (
            .O(N__31381),
            .I(N__31374));
    Span4Mux_h I__5919 (
            .O(N__31374),
            .I(N__31368));
    InMux I__5918 (
            .O(N__31373),
            .I(N__31363));
    InMux I__5917 (
            .O(N__31372),
            .I(N__31363));
    InMux I__5916 (
            .O(N__31371),
            .I(N__31360));
    Odrv4 I__5915 (
            .O(N__31368),
            .I(\current_shift_inst.S1_riseZ0 ));
    LocalMux I__5914 (
            .O(N__31363),
            .I(\current_shift_inst.S1_riseZ0 ));
    LocalMux I__5913 (
            .O(N__31360),
            .I(\current_shift_inst.S1_riseZ0 ));
    InMux I__5912 (
            .O(N__31353),
            .I(N__31350));
    LocalMux I__5911 (
            .O(N__31350),
            .I(N__31347));
    Odrv4 I__5910 (
            .O(N__31347),
            .I(\current_shift_inst.N_199 ));
    CascadeMux I__5909 (
            .O(N__31344),
            .I(N__31339));
    CascadeMux I__5908 (
            .O(N__31343),
            .I(N__31336));
    InMux I__5907 (
            .O(N__31342),
            .I(N__31328));
    InMux I__5906 (
            .O(N__31339),
            .I(N__31328));
    InMux I__5905 (
            .O(N__31336),
            .I(N__31323));
    InMux I__5904 (
            .O(N__31335),
            .I(N__31323));
    InMux I__5903 (
            .O(N__31334),
            .I(N__31317));
    InMux I__5902 (
            .O(N__31333),
            .I(N__31317));
    LocalMux I__5901 (
            .O(N__31328),
            .I(N__31312));
    LocalMux I__5900 (
            .O(N__31323),
            .I(N__31312));
    InMux I__5899 (
            .O(N__31322),
            .I(N__31309));
    LocalMux I__5898 (
            .O(N__31317),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    Odrv4 I__5897 (
            .O(N__31312),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__5896 (
            .O(N__31309),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    InMux I__5895 (
            .O(N__31302),
            .I(N__31298));
    InMux I__5894 (
            .O(N__31301),
            .I(N__31295));
    LocalMux I__5893 (
            .O(N__31298),
            .I(measured_delay_hc_28));
    LocalMux I__5892 (
            .O(N__31295),
            .I(measured_delay_hc_28));
    CascadeMux I__5891 (
            .O(N__31290),
            .I(N__31287));
    InMux I__5890 (
            .O(N__31287),
            .I(N__31283));
    InMux I__5889 (
            .O(N__31286),
            .I(N__31280));
    LocalMux I__5888 (
            .O(N__31283),
            .I(measured_delay_hc_29));
    LocalMux I__5887 (
            .O(N__31280),
            .I(measured_delay_hc_29));
    CascadeMux I__5886 (
            .O(N__31275),
            .I(N__31271));
    InMux I__5885 (
            .O(N__31274),
            .I(N__31268));
    InMux I__5884 (
            .O(N__31271),
            .I(N__31265));
    LocalMux I__5883 (
            .O(N__31268),
            .I(measured_delay_hc_30));
    LocalMux I__5882 (
            .O(N__31265),
            .I(measured_delay_hc_30));
    InMux I__5881 (
            .O(N__31260),
            .I(N__31257));
    LocalMux I__5880 (
            .O(N__31257),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ));
    CascadeMux I__5879 (
            .O(N__31254),
            .I(N__31251));
    InMux I__5878 (
            .O(N__31251),
            .I(N__31248));
    LocalMux I__5877 (
            .O(N__31248),
            .I(N__31245));
    Odrv12 I__5876 (
            .O(N__31245),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    InMux I__5875 (
            .O(N__31242),
            .I(N__31239));
    LocalMux I__5874 (
            .O(N__31239),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    CascadeMux I__5873 (
            .O(N__31236),
            .I(N__31233));
    InMux I__5872 (
            .O(N__31233),
            .I(N__31230));
    LocalMux I__5871 (
            .O(N__31230),
            .I(N__31227));
    Span4Mux_v I__5870 (
            .O(N__31227),
            .I(N__31224));
    Odrv4 I__5869 (
            .O(N__31224),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__5868 (
            .O(N__31221),
            .I(N__31218));
    LocalMux I__5867 (
            .O(N__31218),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__5866 (
            .O(N__31215),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__5865 (
            .O(N__31212),
            .I(N__31209));
    LocalMux I__5864 (
            .O(N__31209),
            .I(N__31206));
    Odrv4 I__5863 (
            .O(N__31206),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10 ));
    InMux I__5862 (
            .O(N__31203),
            .I(N__31200));
    LocalMux I__5861 (
            .O(N__31200),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ));
    InMux I__5860 (
            .O(N__31197),
            .I(N__31194));
    LocalMux I__5859 (
            .O(N__31194),
            .I(\current_shift_inst.S3_sync_prevZ0 ));
    InMux I__5858 (
            .O(N__31191),
            .I(N__31187));
    CascadeMux I__5857 (
            .O(N__31190),
            .I(N__31184));
    LocalMux I__5856 (
            .O(N__31187),
            .I(N__31181));
    InMux I__5855 (
            .O(N__31184),
            .I(N__31178));
    Odrv4 I__5854 (
            .O(N__31181),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    LocalMux I__5853 (
            .O(N__31178),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    CascadeMux I__5852 (
            .O(N__31173),
            .I(N__31170));
    InMux I__5851 (
            .O(N__31170),
            .I(N__31167));
    LocalMux I__5850 (
            .O(N__31167),
            .I(N__31164));
    Odrv4 I__5849 (
            .O(N__31164),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__5848 (
            .O(N__31161),
            .I(N__31158));
    LocalMux I__5847 (
            .O(N__31158),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__5846 (
            .O(N__31155),
            .I(N__31152));
    InMux I__5845 (
            .O(N__31152),
            .I(N__31149));
    LocalMux I__5844 (
            .O(N__31149),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__5843 (
            .O(N__31146),
            .I(N__31143));
    LocalMux I__5842 (
            .O(N__31143),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__5841 (
            .O(N__31140),
            .I(N__31137));
    InMux I__5840 (
            .O(N__31137),
            .I(N__31134));
    LocalMux I__5839 (
            .O(N__31134),
            .I(N__31131));
    Odrv4 I__5838 (
            .O(N__31131),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__5837 (
            .O(N__31128),
            .I(N__31125));
    LocalMux I__5836 (
            .O(N__31125),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__5835 (
            .O(N__31122),
            .I(N__31119));
    InMux I__5834 (
            .O(N__31119),
            .I(N__31116));
    LocalMux I__5833 (
            .O(N__31116),
            .I(N__31113));
    Span4Mux_h I__5832 (
            .O(N__31113),
            .I(N__31110));
    Odrv4 I__5831 (
            .O(N__31110),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__5830 (
            .O(N__31107),
            .I(N__31104));
    LocalMux I__5829 (
            .O(N__31104),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__5828 (
            .O(N__31101),
            .I(N__31098));
    InMux I__5827 (
            .O(N__31098),
            .I(N__31095));
    LocalMux I__5826 (
            .O(N__31095),
            .I(N__31092));
    Odrv4 I__5825 (
            .O(N__31092),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__5824 (
            .O(N__31089),
            .I(N__31086));
    LocalMux I__5823 (
            .O(N__31086),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__5822 (
            .O(N__31083),
            .I(N__31080));
    InMux I__5821 (
            .O(N__31080),
            .I(N__31077));
    LocalMux I__5820 (
            .O(N__31077),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__5819 (
            .O(N__31074),
            .I(N__31071));
    LocalMux I__5818 (
            .O(N__31071),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__5817 (
            .O(N__31068),
            .I(N__31065));
    InMux I__5816 (
            .O(N__31065),
            .I(N__31062));
    LocalMux I__5815 (
            .O(N__31062),
            .I(N__31059));
    Odrv4 I__5814 (
            .O(N__31059),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__5813 (
            .O(N__31056),
            .I(N__31053));
    LocalMux I__5812 (
            .O(N__31053),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    CascadeMux I__5811 (
            .O(N__31050),
            .I(N__31047));
    InMux I__5810 (
            .O(N__31047),
            .I(N__31044));
    LocalMux I__5809 (
            .O(N__31044),
            .I(N__31041));
    Odrv4 I__5808 (
            .O(N__31041),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__5807 (
            .O(N__31038),
            .I(N__31035));
    LocalMux I__5806 (
            .O(N__31035),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__5805 (
            .O(N__31032),
            .I(N__31029));
    InMux I__5804 (
            .O(N__31029),
            .I(N__31026));
    LocalMux I__5803 (
            .O(N__31026),
            .I(N__31023));
    Odrv4 I__5802 (
            .O(N__31023),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__5801 (
            .O(N__31020),
            .I(N__31017));
    LocalMux I__5800 (
            .O(N__31017),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__5799 (
            .O(N__31014),
            .I(N__31011));
    InMux I__5798 (
            .O(N__31011),
            .I(N__31008));
    LocalMux I__5797 (
            .O(N__31008),
            .I(N__31005));
    Span4Mux_h I__5796 (
            .O(N__31005),
            .I(N__31002));
    Odrv4 I__5795 (
            .O(N__31002),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__5794 (
            .O(N__30999),
            .I(N__30996));
    LocalMux I__5793 (
            .O(N__30996),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__5792 (
            .O(N__30993),
            .I(N__30990));
    InMux I__5791 (
            .O(N__30990),
            .I(N__30987));
    LocalMux I__5790 (
            .O(N__30987),
            .I(N__30984));
    Span4Mux_v I__5789 (
            .O(N__30984),
            .I(N__30981));
    Odrv4 I__5788 (
            .O(N__30981),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ));
    InMux I__5787 (
            .O(N__30978),
            .I(N__30975));
    LocalMux I__5786 (
            .O(N__30975),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__5785 (
            .O(N__30972),
            .I(N__30969));
    InMux I__5784 (
            .O(N__30969),
            .I(N__30966));
    LocalMux I__5783 (
            .O(N__30966),
            .I(N__30963));
    Odrv4 I__5782 (
            .O(N__30963),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__5781 (
            .O(N__30960),
            .I(N__30957));
    LocalMux I__5780 (
            .O(N__30957),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__5779 (
            .O(N__30954),
            .I(N__30951));
    InMux I__5778 (
            .O(N__30951),
            .I(N__30948));
    LocalMux I__5777 (
            .O(N__30948),
            .I(N__30945));
    Span4Mux_v I__5776 (
            .O(N__30945),
            .I(N__30942));
    Odrv4 I__5775 (
            .O(N__30942),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    InMux I__5774 (
            .O(N__30939),
            .I(N__30936));
    LocalMux I__5773 (
            .O(N__30936),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__5772 (
            .O(N__30933),
            .I(N__30930));
    InMux I__5771 (
            .O(N__30930),
            .I(N__30927));
    LocalMux I__5770 (
            .O(N__30927),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__5769 (
            .O(N__30924),
            .I(N__30921));
    LocalMux I__5768 (
            .O(N__30921),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__5767 (
            .O(N__30918),
            .I(N__30915));
    InMux I__5766 (
            .O(N__30915),
            .I(N__30912));
    LocalMux I__5765 (
            .O(N__30912),
            .I(N__30909));
    Odrv4 I__5764 (
            .O(N__30909),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__5763 (
            .O(N__30906),
            .I(N__30903));
    LocalMux I__5762 (
            .O(N__30903),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__5761 (
            .O(N__30900),
            .I(N__30897));
    LocalMux I__5760 (
            .O(N__30897),
            .I(N__30894));
    Odrv12 I__5759 (
            .O(N__30894),
            .I(il_max_comp1_D1));
    CascadeMux I__5758 (
            .O(N__30891),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_ ));
    CEMux I__5757 (
            .O(N__30888),
            .I(N__30878));
    CEMux I__5756 (
            .O(N__30887),
            .I(N__30875));
    CEMux I__5755 (
            .O(N__30886),
            .I(N__30872));
    CEMux I__5754 (
            .O(N__30885),
            .I(N__30869));
    CEMux I__5753 (
            .O(N__30884),
            .I(N__30866));
    CEMux I__5752 (
            .O(N__30883),
            .I(N__30863));
    CEMux I__5751 (
            .O(N__30882),
            .I(N__30860));
    CEMux I__5750 (
            .O(N__30881),
            .I(N__30857));
    LocalMux I__5749 (
            .O(N__30878),
            .I(N__30853));
    LocalMux I__5748 (
            .O(N__30875),
            .I(N__30850));
    LocalMux I__5747 (
            .O(N__30872),
            .I(N__30847));
    LocalMux I__5746 (
            .O(N__30869),
            .I(N__30844));
    LocalMux I__5745 (
            .O(N__30866),
            .I(N__30841));
    LocalMux I__5744 (
            .O(N__30863),
            .I(N__30838));
    LocalMux I__5743 (
            .O(N__30860),
            .I(N__30835));
    LocalMux I__5742 (
            .O(N__30857),
            .I(N__30832));
    CEMux I__5741 (
            .O(N__30856),
            .I(N__30829));
    Span12Mux_s10_h I__5740 (
            .O(N__30853),
            .I(N__30826));
    Span4Mux_v I__5739 (
            .O(N__30850),
            .I(N__30823));
    Span4Mux_v I__5738 (
            .O(N__30847),
            .I(N__30818));
    Span4Mux_v I__5737 (
            .O(N__30844),
            .I(N__30818));
    Span4Mux_v I__5736 (
            .O(N__30841),
            .I(N__30811));
    Span4Mux_h I__5735 (
            .O(N__30838),
            .I(N__30811));
    Span4Mux_v I__5734 (
            .O(N__30835),
            .I(N__30811));
    Span4Mux_v I__5733 (
            .O(N__30832),
            .I(N__30806));
    LocalMux I__5732 (
            .O(N__30829),
            .I(N__30806));
    Odrv12 I__5731 (
            .O(N__30826),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5730 (
            .O(N__30823),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5729 (
            .O(N__30818),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5728 (
            .O(N__30811),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5727 (
            .O(N__30806),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__5726 (
            .O(N__30795),
            .I(N__30792));
    LocalMux I__5725 (
            .O(N__30792),
            .I(N__30789));
    Odrv4 I__5724 (
            .O(N__30789),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__5723 (
            .O(N__30786),
            .I(N__30783));
    InMux I__5722 (
            .O(N__30783),
            .I(N__30780));
    LocalMux I__5721 (
            .O(N__30780),
            .I(N__30777));
    Odrv4 I__5720 (
            .O(N__30777),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__5719 (
            .O(N__30774),
            .I(N__30771));
    LocalMux I__5718 (
            .O(N__30771),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__5717 (
            .O(N__30768),
            .I(N__30765));
    InMux I__5716 (
            .O(N__30765),
            .I(N__30762));
    LocalMux I__5715 (
            .O(N__30762),
            .I(N__30759));
    Span4Mux_v I__5714 (
            .O(N__30759),
            .I(N__30756));
    Sp12to4 I__5713 (
            .O(N__30756),
            .I(N__30753));
    Odrv12 I__5712 (
            .O(N__30753),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__5711 (
            .O(N__30750),
            .I(N__30747));
    LocalMux I__5710 (
            .O(N__30747),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__5709 (
            .O(N__30744),
            .I(N__30741));
    InMux I__5708 (
            .O(N__30741),
            .I(N__30738));
    LocalMux I__5707 (
            .O(N__30738),
            .I(N__30735));
    Span4Mux_h I__5706 (
            .O(N__30735),
            .I(N__30732));
    Odrv4 I__5705 (
            .O(N__30732),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ));
    InMux I__5704 (
            .O(N__30729),
            .I(N__30726));
    LocalMux I__5703 (
            .O(N__30726),
            .I(N__30723));
    Span4Mux_h I__5702 (
            .O(N__30723),
            .I(N__30719));
    InMux I__5701 (
            .O(N__30722),
            .I(N__30716));
    Span4Mux_v I__5700 (
            .O(N__30719),
            .I(N__30713));
    LocalMux I__5699 (
            .O(N__30716),
            .I(\current_shift_inst.z_31 ));
    Odrv4 I__5698 (
            .O(N__30713),
            .I(\current_shift_inst.z_31 ));
    CascadeMux I__5697 (
            .O(N__30708),
            .I(N__30704));
    InMux I__5696 (
            .O(N__30707),
            .I(N__30701));
    InMux I__5695 (
            .O(N__30704),
            .I(N__30698));
    LocalMux I__5694 (
            .O(N__30701),
            .I(N__30693));
    LocalMux I__5693 (
            .O(N__30698),
            .I(N__30693));
    Span4Mux_h I__5692 (
            .O(N__30693),
            .I(N__30690));
    Span4Mux_v I__5691 (
            .O(N__30690),
            .I(N__30687));
    Odrv4 I__5690 (
            .O(N__30687),
            .I(\current_shift_inst.z_i_31 ));
    CascadeMux I__5689 (
            .O(N__30684),
            .I(N__30680));
    InMux I__5688 (
            .O(N__30683),
            .I(N__30676));
    InMux I__5687 (
            .O(N__30680),
            .I(N__30671));
    InMux I__5686 (
            .O(N__30679),
            .I(N__30671));
    LocalMux I__5685 (
            .O(N__30676),
            .I(N__30668));
    LocalMux I__5684 (
            .O(N__30671),
            .I(N__30665));
    Span12Mux_s11_v I__5683 (
            .O(N__30668),
            .I(N__30661));
    Span4Mux_v I__5682 (
            .O(N__30665),
            .I(N__30658));
    InMux I__5681 (
            .O(N__30664),
            .I(N__30655));
    Odrv12 I__5680 (
            .O(N__30661),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    Odrv4 I__5679 (
            .O(N__30658),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    LocalMux I__5678 (
            .O(N__30655),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    CascadeMux I__5677 (
            .O(N__30648),
            .I(N__30642));
    CascadeMux I__5676 (
            .O(N__30647),
            .I(N__30639));
    InMux I__5675 (
            .O(N__30646),
            .I(N__30636));
    InMux I__5674 (
            .O(N__30645),
            .I(N__30631));
    InMux I__5673 (
            .O(N__30642),
            .I(N__30631));
    InMux I__5672 (
            .O(N__30639),
            .I(N__30628));
    LocalMux I__5671 (
            .O(N__30636),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    LocalMux I__5670 (
            .O(N__30631),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    LocalMux I__5669 (
            .O(N__30628),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    InMux I__5668 (
            .O(N__30621),
            .I(N__30618));
    LocalMux I__5667 (
            .O(N__30618),
            .I(N__30615));
    Span4Mux_h I__5666 (
            .O(N__30615),
            .I(N__30612));
    Odrv4 I__5665 (
            .O(N__30612),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ));
    CascadeMux I__5664 (
            .O(N__30609),
            .I(N__30606));
    InMux I__5663 (
            .O(N__30606),
            .I(N__30603));
    LocalMux I__5662 (
            .O(N__30603),
            .I(N__30600));
    Span4Mux_h I__5661 (
            .O(N__30600),
            .I(N__30597));
    Odrv4 I__5660 (
            .O(N__30597),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ));
    InMux I__5659 (
            .O(N__30594),
            .I(N__30589));
    InMux I__5658 (
            .O(N__30593),
            .I(N__30586));
    CascadeMux I__5657 (
            .O(N__30592),
            .I(N__30582));
    LocalMux I__5656 (
            .O(N__30589),
            .I(N__30574));
    LocalMux I__5655 (
            .O(N__30586),
            .I(N__30574));
    InMux I__5654 (
            .O(N__30585),
            .I(N__30571));
    InMux I__5653 (
            .O(N__30582),
            .I(N__30568));
    InMux I__5652 (
            .O(N__30581),
            .I(N__30565));
    CascadeMux I__5651 (
            .O(N__30580),
            .I(N__30561));
    CascadeMux I__5650 (
            .O(N__30579),
            .I(N__30557));
    Span4Mux_v I__5649 (
            .O(N__30574),
            .I(N__30552));
    LocalMux I__5648 (
            .O(N__30571),
            .I(N__30552));
    LocalMux I__5647 (
            .O(N__30568),
            .I(N__30549));
    LocalMux I__5646 (
            .O(N__30565),
            .I(N__30546));
    InMux I__5645 (
            .O(N__30564),
            .I(N__30537));
    InMux I__5644 (
            .O(N__30561),
            .I(N__30537));
    InMux I__5643 (
            .O(N__30560),
            .I(N__30537));
    InMux I__5642 (
            .O(N__30557),
            .I(N__30537));
    Span4Mux_v I__5641 (
            .O(N__30552),
            .I(N__30534));
    Odrv4 I__5640 (
            .O(N__30549),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5639 (
            .O(N__30546),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__5638 (
            .O(N__30537),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5637 (
            .O(N__30534),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__5636 (
            .O(N__30525),
            .I(N__30521));
    InMux I__5635 (
            .O(N__30524),
            .I(N__30518));
    LocalMux I__5634 (
            .O(N__30521),
            .I(N__30514));
    LocalMux I__5633 (
            .O(N__30518),
            .I(N__30511));
    InMux I__5632 (
            .O(N__30517),
            .I(N__30508));
    Odrv4 I__5631 (
            .O(N__30514),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    Odrv4 I__5630 (
            .O(N__30511),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    LocalMux I__5629 (
            .O(N__30508),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    CascadeMux I__5628 (
            .O(N__30501),
            .I(N__30497));
    CascadeMux I__5627 (
            .O(N__30500),
            .I(N__30494));
    InMux I__5626 (
            .O(N__30497),
            .I(N__30491));
    InMux I__5625 (
            .O(N__30494),
            .I(N__30488));
    LocalMux I__5624 (
            .O(N__30491),
            .I(N__30483));
    LocalMux I__5623 (
            .O(N__30488),
            .I(N__30483));
    Span4Mux_h I__5622 (
            .O(N__30483),
            .I(N__30480));
    Odrv4 I__5621 (
            .O(N__30480),
            .I(\current_shift_inst.elapsed_time_ns_phase_31 ));
    InMux I__5620 (
            .O(N__30477),
            .I(N__30474));
    LocalMux I__5619 (
            .O(N__30474),
            .I(N__30470));
    InMux I__5618 (
            .O(N__30473),
            .I(N__30466));
    Span4Mux_h I__5617 (
            .O(N__30470),
            .I(N__30463));
    InMux I__5616 (
            .O(N__30469),
            .I(N__30460));
    LocalMux I__5615 (
            .O(N__30466),
            .I(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ));
    Odrv4 I__5614 (
            .O(N__30463),
            .I(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ));
    LocalMux I__5613 (
            .O(N__30460),
            .I(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ));
    InMux I__5612 (
            .O(N__30453),
            .I(N__30450));
    LocalMux I__5611 (
            .O(N__30450),
            .I(N__30447));
    Span4Mux_v I__5610 (
            .O(N__30447),
            .I(N__30444));
    Odrv4 I__5609 (
            .O(N__30444),
            .I(\current_shift_inst.un38_control_input_0_axb_31 ));
    InMux I__5608 (
            .O(N__30441),
            .I(N__30436));
    InMux I__5607 (
            .O(N__30440),
            .I(N__30433));
    InMux I__5606 (
            .O(N__30439),
            .I(N__30429));
    LocalMux I__5605 (
            .O(N__30436),
            .I(N__30426));
    LocalMux I__5604 (
            .O(N__30433),
            .I(N__30423));
    InMux I__5603 (
            .O(N__30432),
            .I(N__30420));
    LocalMux I__5602 (
            .O(N__30429),
            .I(N__30417));
    Span4Mux_h I__5601 (
            .O(N__30426),
            .I(N__30412));
    Span4Mux_h I__5600 (
            .O(N__30423),
            .I(N__30412));
    LocalMux I__5599 (
            .O(N__30420),
            .I(N__30409));
    Odrv12 I__5598 (
            .O(N__30417),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    Odrv4 I__5597 (
            .O(N__30412),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    Odrv4 I__5596 (
            .O(N__30409),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    InMux I__5595 (
            .O(N__30402),
            .I(N__30399));
    LocalMux I__5594 (
            .O(N__30399),
            .I(N__30395));
    CascadeMux I__5593 (
            .O(N__30398),
            .I(N__30390));
    Span4Mux_h I__5592 (
            .O(N__30395),
            .I(N__30387));
    InMux I__5591 (
            .O(N__30394),
            .I(N__30384));
    InMux I__5590 (
            .O(N__30393),
            .I(N__30381));
    InMux I__5589 (
            .O(N__30390),
            .I(N__30378));
    Odrv4 I__5588 (
            .O(N__30387),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    LocalMux I__5587 (
            .O(N__30384),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    LocalMux I__5586 (
            .O(N__30381),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    LocalMux I__5585 (
            .O(N__30378),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    CascadeMux I__5584 (
            .O(N__30369),
            .I(N__30366));
    InMux I__5583 (
            .O(N__30366),
            .I(N__30363));
    LocalMux I__5582 (
            .O(N__30363),
            .I(N__30360));
    Span4Mux_h I__5581 (
            .O(N__30360),
            .I(N__30357));
    Span4Mux_v I__5580 (
            .O(N__30357),
            .I(N__30354));
    Odrv4 I__5579 (
            .O(N__30354),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ));
    CascadeMux I__5578 (
            .O(N__30351),
            .I(N__30347));
    InMux I__5577 (
            .O(N__30350),
            .I(N__30343));
    InMux I__5576 (
            .O(N__30347),
            .I(N__30338));
    InMux I__5575 (
            .O(N__30346),
            .I(N__30338));
    LocalMux I__5574 (
            .O(N__30343),
            .I(N__30335));
    LocalMux I__5573 (
            .O(N__30338),
            .I(N__30332));
    Span4Mux_v I__5572 (
            .O(N__30335),
            .I(N__30328));
    Span4Mux_h I__5571 (
            .O(N__30332),
            .I(N__30325));
    InMux I__5570 (
            .O(N__30331),
            .I(N__30322));
    Odrv4 I__5569 (
            .O(N__30328),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    Odrv4 I__5568 (
            .O(N__30325),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    LocalMux I__5567 (
            .O(N__30322),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    InMux I__5566 (
            .O(N__30315),
            .I(N__30305));
    InMux I__5565 (
            .O(N__30314),
            .I(N__30305));
    InMux I__5564 (
            .O(N__30313),
            .I(N__30305));
    CascadeMux I__5563 (
            .O(N__30312),
            .I(N__30302));
    LocalMux I__5562 (
            .O(N__30305),
            .I(N__30299));
    InMux I__5561 (
            .O(N__30302),
            .I(N__30296));
    Odrv4 I__5560 (
            .O(N__30299),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    LocalMux I__5559 (
            .O(N__30296),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    CascadeMux I__5558 (
            .O(N__30291),
            .I(N__30286));
    InMux I__5557 (
            .O(N__30290),
            .I(N__30281));
    InMux I__5556 (
            .O(N__30289),
            .I(N__30281));
    InMux I__5555 (
            .O(N__30286),
            .I(N__30277));
    LocalMux I__5554 (
            .O(N__30281),
            .I(N__30274));
    CascadeMux I__5553 (
            .O(N__30280),
            .I(N__30271));
    LocalMux I__5552 (
            .O(N__30277),
            .I(N__30268));
    Span4Mux_h I__5551 (
            .O(N__30274),
            .I(N__30265));
    InMux I__5550 (
            .O(N__30271),
            .I(N__30262));
    Odrv4 I__5549 (
            .O(N__30268),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    Odrv4 I__5548 (
            .O(N__30265),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    LocalMux I__5547 (
            .O(N__30262),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    CascadeMux I__5546 (
            .O(N__30255),
            .I(N__30251));
    InMux I__5545 (
            .O(N__30254),
            .I(N__30243));
    InMux I__5544 (
            .O(N__30251),
            .I(N__30243));
    InMux I__5543 (
            .O(N__30250),
            .I(N__30243));
    LocalMux I__5542 (
            .O(N__30243),
            .I(N__30240));
    Span4Mux_v I__5541 (
            .O(N__30240),
            .I(N__30236));
    InMux I__5540 (
            .O(N__30239),
            .I(N__30233));
    Odrv4 I__5539 (
            .O(N__30236),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    LocalMux I__5538 (
            .O(N__30233),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    InMux I__5537 (
            .O(N__30228),
            .I(N__30225));
    LocalMux I__5536 (
            .O(N__30225),
            .I(N__30222));
    Span4Mux_h I__5535 (
            .O(N__30222),
            .I(N__30219));
    Span4Mux_v I__5534 (
            .O(N__30219),
            .I(N__30216));
    Odrv4 I__5533 (
            .O(N__30216),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ));
    InMux I__5532 (
            .O(N__30213),
            .I(bfn_11_19_0_));
    InMux I__5531 (
            .O(N__30210),
            .I(\current_shift_inst.un4_control_input_cry_25 ));
    InMux I__5530 (
            .O(N__30207),
            .I(\current_shift_inst.un4_control_input_cry_26 ));
    CascadeMux I__5529 (
            .O(N__30204),
            .I(N__30200));
    CascadeMux I__5528 (
            .O(N__30203),
            .I(N__30197));
    InMux I__5527 (
            .O(N__30200),
            .I(N__30189));
    InMux I__5526 (
            .O(N__30197),
            .I(N__30189));
    InMux I__5525 (
            .O(N__30196),
            .I(N__30189));
    LocalMux I__5524 (
            .O(N__30189),
            .I(N__30185));
    CascadeMux I__5523 (
            .O(N__30188),
            .I(N__30182));
    Span4Mux_h I__5522 (
            .O(N__30185),
            .I(N__30179));
    InMux I__5521 (
            .O(N__30182),
            .I(N__30176));
    Odrv4 I__5520 (
            .O(N__30179),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    LocalMux I__5519 (
            .O(N__30176),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    InMux I__5518 (
            .O(N__30171),
            .I(\current_shift_inst.un4_control_input_cry_27 ));
    InMux I__5517 (
            .O(N__30168),
            .I(N__30159));
    InMux I__5516 (
            .O(N__30167),
            .I(N__30159));
    InMux I__5515 (
            .O(N__30166),
            .I(N__30159));
    LocalMux I__5514 (
            .O(N__30159),
            .I(N__30155));
    CascadeMux I__5513 (
            .O(N__30158),
            .I(N__30152));
    Span4Mux_v I__5512 (
            .O(N__30155),
            .I(N__30149));
    InMux I__5511 (
            .O(N__30152),
            .I(N__30146));
    Odrv4 I__5510 (
            .O(N__30149),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    LocalMux I__5509 (
            .O(N__30146),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    InMux I__5508 (
            .O(N__30141),
            .I(\current_shift_inst.un4_control_input_cry_28 ));
    InMux I__5507 (
            .O(N__30138),
            .I(N__30132));
    InMux I__5506 (
            .O(N__30137),
            .I(N__30132));
    LocalMux I__5505 (
            .O(N__30132),
            .I(N__30129));
    Span4Mux_v I__5504 (
            .O(N__30129),
            .I(N__30125));
    InMux I__5503 (
            .O(N__30128),
            .I(N__30122));
    Odrv4 I__5502 (
            .O(N__30125),
            .I(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ));
    LocalMux I__5501 (
            .O(N__30122),
            .I(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ));
    InMux I__5500 (
            .O(N__30117),
            .I(\current_shift_inst.un4_control_input_cry_29 ));
    InMux I__5499 (
            .O(N__30114),
            .I(\current_shift_inst.un4_control_input_cry_30 ));
    InMux I__5498 (
            .O(N__30111),
            .I(N__30108));
    LocalMux I__5497 (
            .O(N__30108),
            .I(N__30105));
    Span4Mux_h I__5496 (
            .O(N__30105),
            .I(N__30102));
    Odrv4 I__5495 (
            .O(N__30102),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ));
    InMux I__5494 (
            .O(N__30099),
            .I(N__30095));
    InMux I__5493 (
            .O(N__30098),
            .I(N__30090));
    LocalMux I__5492 (
            .O(N__30095),
            .I(N__30087));
    InMux I__5491 (
            .O(N__30094),
            .I(N__30084));
    InMux I__5490 (
            .O(N__30093),
            .I(N__30081));
    LocalMux I__5489 (
            .O(N__30090),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    Odrv12 I__5488 (
            .O(N__30087),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    LocalMux I__5487 (
            .O(N__30084),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    LocalMux I__5486 (
            .O(N__30081),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    InMux I__5485 (
            .O(N__30072),
            .I(N__30067));
    CascadeMux I__5484 (
            .O(N__30071),
            .I(N__30064));
    InMux I__5483 (
            .O(N__30070),
            .I(N__30061));
    LocalMux I__5482 (
            .O(N__30067),
            .I(N__30058));
    InMux I__5481 (
            .O(N__30064),
            .I(N__30054));
    LocalMux I__5480 (
            .O(N__30061),
            .I(N__30051));
    Span4Mux_h I__5479 (
            .O(N__30058),
            .I(N__30048));
    InMux I__5478 (
            .O(N__30057),
            .I(N__30045));
    LocalMux I__5477 (
            .O(N__30054),
            .I(N__30042));
    Span4Mux_h I__5476 (
            .O(N__30051),
            .I(N__30037));
    Span4Mux_v I__5475 (
            .O(N__30048),
            .I(N__30037));
    LocalMux I__5474 (
            .O(N__30045),
            .I(N__30034));
    Odrv12 I__5473 (
            .O(N__30042),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    Odrv4 I__5472 (
            .O(N__30037),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    Odrv4 I__5471 (
            .O(N__30034),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    InMux I__5470 (
            .O(N__30027),
            .I(N__30024));
    LocalMux I__5469 (
            .O(N__30024),
            .I(N__30021));
    Span4Mux_h I__5468 (
            .O(N__30021),
            .I(N__30018));
    Odrv4 I__5467 (
            .O(N__30018),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ));
    CascadeMux I__5466 (
            .O(N__30015),
            .I(N__30012));
    InMux I__5465 (
            .O(N__30012),
            .I(N__30003));
    InMux I__5464 (
            .O(N__30011),
            .I(N__30003));
    InMux I__5463 (
            .O(N__30010),
            .I(N__30003));
    LocalMux I__5462 (
            .O(N__30003),
            .I(N__29999));
    CascadeMux I__5461 (
            .O(N__30002),
            .I(N__29996));
    Span4Mux_h I__5460 (
            .O(N__29999),
            .I(N__29993));
    InMux I__5459 (
            .O(N__29996),
            .I(N__29990));
    Odrv4 I__5458 (
            .O(N__29993),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    LocalMux I__5457 (
            .O(N__29990),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    InMux I__5456 (
            .O(N__29985),
            .I(\current_shift_inst.un4_control_input_cry_15 ));
    CascadeMux I__5455 (
            .O(N__29982),
            .I(N__29979));
    InMux I__5454 (
            .O(N__29979),
            .I(N__29970));
    InMux I__5453 (
            .O(N__29978),
            .I(N__29970));
    InMux I__5452 (
            .O(N__29977),
            .I(N__29970));
    LocalMux I__5451 (
            .O(N__29970),
            .I(N__29966));
    CascadeMux I__5450 (
            .O(N__29969),
            .I(N__29963));
    Span4Mux_h I__5449 (
            .O(N__29966),
            .I(N__29960));
    InMux I__5448 (
            .O(N__29963),
            .I(N__29957));
    Odrv4 I__5447 (
            .O(N__29960),
            .I(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ));
    LocalMux I__5446 (
            .O(N__29957),
            .I(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ));
    InMux I__5445 (
            .O(N__29952),
            .I(bfn_11_18_0_));
    CascadeMux I__5444 (
            .O(N__29949),
            .I(N__29946));
    InMux I__5443 (
            .O(N__29946),
            .I(N__29943));
    LocalMux I__5442 (
            .O(N__29943),
            .I(N__29938));
    InMux I__5441 (
            .O(N__29942),
            .I(N__29935));
    InMux I__5440 (
            .O(N__29941),
            .I(N__29932));
    Span4Mux_v I__5439 (
            .O(N__29938),
            .I(N__29924));
    LocalMux I__5438 (
            .O(N__29935),
            .I(N__29924));
    LocalMux I__5437 (
            .O(N__29932),
            .I(N__29924));
    CascadeMux I__5436 (
            .O(N__29931),
            .I(N__29921));
    Span4Mux_h I__5435 (
            .O(N__29924),
            .I(N__29918));
    InMux I__5434 (
            .O(N__29921),
            .I(N__29915));
    Odrv4 I__5433 (
            .O(N__29918),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    LocalMux I__5432 (
            .O(N__29915),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    InMux I__5431 (
            .O(N__29910),
            .I(\current_shift_inst.un4_control_input_cry_17 ));
    CascadeMux I__5430 (
            .O(N__29907),
            .I(N__29904));
    InMux I__5429 (
            .O(N__29904),
            .I(N__29899));
    InMux I__5428 (
            .O(N__29903),
            .I(N__29894));
    InMux I__5427 (
            .O(N__29902),
            .I(N__29894));
    LocalMux I__5426 (
            .O(N__29899),
            .I(N__29890));
    LocalMux I__5425 (
            .O(N__29894),
            .I(N__29887));
    CascadeMux I__5424 (
            .O(N__29893),
            .I(N__29884));
    Span4Mux_h I__5423 (
            .O(N__29890),
            .I(N__29881));
    Span4Mux_v I__5422 (
            .O(N__29887),
            .I(N__29878));
    InMux I__5421 (
            .O(N__29884),
            .I(N__29875));
    Odrv4 I__5420 (
            .O(N__29881),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    Odrv4 I__5419 (
            .O(N__29878),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    LocalMux I__5418 (
            .O(N__29875),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    InMux I__5417 (
            .O(N__29868),
            .I(\current_shift_inst.un4_control_input_cry_18 ));
    CascadeMux I__5416 (
            .O(N__29865),
            .I(N__29862));
    InMux I__5415 (
            .O(N__29862),
            .I(N__29853));
    InMux I__5414 (
            .O(N__29861),
            .I(N__29853));
    InMux I__5413 (
            .O(N__29860),
            .I(N__29853));
    LocalMux I__5412 (
            .O(N__29853),
            .I(N__29849));
    CascadeMux I__5411 (
            .O(N__29852),
            .I(N__29846));
    Span4Mux_h I__5410 (
            .O(N__29849),
            .I(N__29843));
    InMux I__5409 (
            .O(N__29846),
            .I(N__29840));
    Odrv4 I__5408 (
            .O(N__29843),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    LocalMux I__5407 (
            .O(N__29840),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    InMux I__5406 (
            .O(N__29835),
            .I(\current_shift_inst.un4_control_input_cry_19 ));
    InMux I__5405 (
            .O(N__29832),
            .I(N__29823));
    InMux I__5404 (
            .O(N__29831),
            .I(N__29823));
    InMux I__5403 (
            .O(N__29830),
            .I(N__29823));
    LocalMux I__5402 (
            .O(N__29823),
            .I(N__29820));
    Span4Mux_v I__5401 (
            .O(N__29820),
            .I(N__29816));
    InMux I__5400 (
            .O(N__29819),
            .I(N__29813));
    Odrv4 I__5399 (
            .O(N__29816),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    LocalMux I__5398 (
            .O(N__29813),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    InMux I__5397 (
            .O(N__29808),
            .I(\current_shift_inst.un4_control_input_cry_20 ));
    CascadeMux I__5396 (
            .O(N__29805),
            .I(N__29802));
    InMux I__5395 (
            .O(N__29802),
            .I(N__29793));
    InMux I__5394 (
            .O(N__29801),
            .I(N__29793));
    InMux I__5393 (
            .O(N__29800),
            .I(N__29793));
    LocalMux I__5392 (
            .O(N__29793),
            .I(N__29789));
    CascadeMux I__5391 (
            .O(N__29792),
            .I(N__29786));
    Span4Mux_v I__5390 (
            .O(N__29789),
            .I(N__29783));
    InMux I__5389 (
            .O(N__29786),
            .I(N__29780));
    Odrv4 I__5388 (
            .O(N__29783),
            .I(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ));
    LocalMux I__5387 (
            .O(N__29780),
            .I(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ));
    InMux I__5386 (
            .O(N__29775),
            .I(\current_shift_inst.un4_control_input_cry_21 ));
    InMux I__5385 (
            .O(N__29772),
            .I(\current_shift_inst.un4_control_input_cry_22 ));
    InMux I__5384 (
            .O(N__29769),
            .I(\current_shift_inst.un4_control_input_cry_23 ));
    InMux I__5383 (
            .O(N__29766),
            .I(N__29763));
    LocalMux I__5382 (
            .O(N__29763),
            .I(\current_shift_inst.un4_control_input_axb_8 ));
    InMux I__5381 (
            .O(N__29760),
            .I(N__29755));
    InMux I__5380 (
            .O(N__29759),
            .I(N__29750));
    InMux I__5379 (
            .O(N__29758),
            .I(N__29750));
    LocalMux I__5378 (
            .O(N__29755),
            .I(N__29744));
    LocalMux I__5377 (
            .O(N__29750),
            .I(N__29744));
    CascadeMux I__5376 (
            .O(N__29749),
            .I(N__29741));
    Span4Mux_h I__5375 (
            .O(N__29744),
            .I(N__29738));
    InMux I__5374 (
            .O(N__29741),
            .I(N__29735));
    Odrv4 I__5373 (
            .O(N__29738),
            .I(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ));
    LocalMux I__5372 (
            .O(N__29735),
            .I(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ));
    InMux I__5371 (
            .O(N__29730),
            .I(\current_shift_inst.un4_control_input_cry_7 ));
    InMux I__5370 (
            .O(N__29727),
            .I(N__29724));
    LocalMux I__5369 (
            .O(N__29724),
            .I(N__29721));
    Odrv4 I__5368 (
            .O(N__29721),
            .I(\current_shift_inst.un4_control_input_axb_9 ));
    CascadeMux I__5367 (
            .O(N__29718),
            .I(N__29714));
    CascadeMux I__5366 (
            .O(N__29717),
            .I(N__29711));
    InMux I__5365 (
            .O(N__29714),
            .I(N__29707));
    InMux I__5364 (
            .O(N__29711),
            .I(N__29702));
    InMux I__5363 (
            .O(N__29710),
            .I(N__29702));
    LocalMux I__5362 (
            .O(N__29707),
            .I(N__29698));
    LocalMux I__5361 (
            .O(N__29702),
            .I(N__29695));
    CascadeMux I__5360 (
            .O(N__29701),
            .I(N__29692));
    Span4Mux_h I__5359 (
            .O(N__29698),
            .I(N__29689));
    Span4Mux_h I__5358 (
            .O(N__29695),
            .I(N__29686));
    InMux I__5357 (
            .O(N__29692),
            .I(N__29683));
    Odrv4 I__5356 (
            .O(N__29689),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    Odrv4 I__5355 (
            .O(N__29686),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    LocalMux I__5354 (
            .O(N__29683),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    InMux I__5353 (
            .O(N__29676),
            .I(bfn_11_17_0_));
    CascadeMux I__5352 (
            .O(N__29673),
            .I(N__29669));
    InMux I__5351 (
            .O(N__29672),
            .I(N__29665));
    InMux I__5350 (
            .O(N__29669),
            .I(N__29660));
    InMux I__5349 (
            .O(N__29668),
            .I(N__29660));
    LocalMux I__5348 (
            .O(N__29665),
            .I(N__29654));
    LocalMux I__5347 (
            .O(N__29660),
            .I(N__29654));
    CascadeMux I__5346 (
            .O(N__29659),
            .I(N__29651));
    Span4Mux_h I__5345 (
            .O(N__29654),
            .I(N__29648));
    InMux I__5344 (
            .O(N__29651),
            .I(N__29645));
    Odrv4 I__5343 (
            .O(N__29648),
            .I(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ));
    LocalMux I__5342 (
            .O(N__29645),
            .I(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ));
    InMux I__5341 (
            .O(N__29640),
            .I(\current_shift_inst.un4_control_input_cry_9 ));
    InMux I__5340 (
            .O(N__29637),
            .I(N__29628));
    InMux I__5339 (
            .O(N__29636),
            .I(N__29628));
    InMux I__5338 (
            .O(N__29635),
            .I(N__29628));
    LocalMux I__5337 (
            .O(N__29628),
            .I(N__29624));
    CascadeMux I__5336 (
            .O(N__29627),
            .I(N__29621));
    Span4Mux_h I__5335 (
            .O(N__29624),
            .I(N__29618));
    InMux I__5334 (
            .O(N__29621),
            .I(N__29615));
    Odrv4 I__5333 (
            .O(N__29618),
            .I(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ));
    LocalMux I__5332 (
            .O(N__29615),
            .I(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ));
    InMux I__5331 (
            .O(N__29610),
            .I(\current_shift_inst.un4_control_input_cry_10 ));
    CascadeMux I__5330 (
            .O(N__29607),
            .I(N__29602));
    InMux I__5329 (
            .O(N__29606),
            .I(N__29599));
    InMux I__5328 (
            .O(N__29605),
            .I(N__29594));
    InMux I__5327 (
            .O(N__29602),
            .I(N__29594));
    LocalMux I__5326 (
            .O(N__29599),
            .I(N__29588));
    LocalMux I__5325 (
            .O(N__29594),
            .I(N__29588));
    CascadeMux I__5324 (
            .O(N__29593),
            .I(N__29585));
    Span4Mux_h I__5323 (
            .O(N__29588),
            .I(N__29582));
    InMux I__5322 (
            .O(N__29585),
            .I(N__29579));
    Odrv4 I__5321 (
            .O(N__29582),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    LocalMux I__5320 (
            .O(N__29579),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    InMux I__5319 (
            .O(N__29574),
            .I(\current_shift_inst.un4_control_input_cry_11 ));
    CascadeMux I__5318 (
            .O(N__29571),
            .I(N__29568));
    InMux I__5317 (
            .O(N__29568),
            .I(N__29564));
    InMux I__5316 (
            .O(N__29567),
            .I(N__29560));
    LocalMux I__5315 (
            .O(N__29564),
            .I(N__29556));
    InMux I__5314 (
            .O(N__29563),
            .I(N__29553));
    LocalMux I__5313 (
            .O(N__29560),
            .I(N__29550));
    CascadeMux I__5312 (
            .O(N__29559),
            .I(N__29547));
    Span4Mux_v I__5311 (
            .O(N__29556),
            .I(N__29540));
    LocalMux I__5310 (
            .O(N__29553),
            .I(N__29540));
    Span4Mux_h I__5309 (
            .O(N__29550),
            .I(N__29540));
    InMux I__5308 (
            .O(N__29547),
            .I(N__29537));
    Odrv4 I__5307 (
            .O(N__29540),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    LocalMux I__5306 (
            .O(N__29537),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    InMux I__5305 (
            .O(N__29532),
            .I(\current_shift_inst.un4_control_input_cry_12 ));
    CascadeMux I__5304 (
            .O(N__29529),
            .I(N__29526));
    InMux I__5303 (
            .O(N__29526),
            .I(N__29523));
    LocalMux I__5302 (
            .O(N__29523),
            .I(N__29518));
    InMux I__5301 (
            .O(N__29522),
            .I(N__29513));
    InMux I__5300 (
            .O(N__29521),
            .I(N__29513));
    Span4Mux_v I__5299 (
            .O(N__29518),
            .I(N__29509));
    LocalMux I__5298 (
            .O(N__29513),
            .I(N__29506));
    CascadeMux I__5297 (
            .O(N__29512),
            .I(N__29503));
    Span4Mux_h I__5296 (
            .O(N__29509),
            .I(N__29498));
    Span4Mux_v I__5295 (
            .O(N__29506),
            .I(N__29498));
    InMux I__5294 (
            .O(N__29503),
            .I(N__29495));
    Odrv4 I__5293 (
            .O(N__29498),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    LocalMux I__5292 (
            .O(N__29495),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    InMux I__5291 (
            .O(N__29490),
            .I(\current_shift_inst.un4_control_input_cry_13 ));
    CascadeMux I__5290 (
            .O(N__29487),
            .I(N__29484));
    InMux I__5289 (
            .O(N__29484),
            .I(N__29477));
    InMux I__5288 (
            .O(N__29483),
            .I(N__29477));
    InMux I__5287 (
            .O(N__29482),
            .I(N__29474));
    LocalMux I__5286 (
            .O(N__29477),
            .I(N__29468));
    LocalMux I__5285 (
            .O(N__29474),
            .I(N__29468));
    CascadeMux I__5284 (
            .O(N__29473),
            .I(N__29465));
    Span4Mux_h I__5283 (
            .O(N__29468),
            .I(N__29462));
    InMux I__5282 (
            .O(N__29465),
            .I(N__29459));
    Odrv4 I__5281 (
            .O(N__29462),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    LocalMux I__5280 (
            .O(N__29459),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    InMux I__5279 (
            .O(N__29454),
            .I(\current_shift_inst.un4_control_input_cry_14 ));
    InMux I__5278 (
            .O(N__29451),
            .I(N__29448));
    LocalMux I__5277 (
            .O(N__29448),
            .I(N__29445));
    Odrv4 I__5276 (
            .O(N__29445),
            .I(\current_shift_inst.un4_control_input_axb_1 ));
    InMux I__5275 (
            .O(N__29442),
            .I(N__29437));
    CascadeMux I__5274 (
            .O(N__29441),
            .I(N__29434));
    InMux I__5273 (
            .O(N__29440),
            .I(N__29431));
    LocalMux I__5272 (
            .O(N__29437),
            .I(N__29428));
    InMux I__5271 (
            .O(N__29434),
            .I(N__29425));
    LocalMux I__5270 (
            .O(N__29431),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    Odrv4 I__5269 (
            .O(N__29428),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    LocalMux I__5268 (
            .O(N__29425),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    CascadeMux I__5267 (
            .O(N__29418),
            .I(N__29415));
    InMux I__5266 (
            .O(N__29415),
            .I(N__29412));
    LocalMux I__5265 (
            .O(N__29412),
            .I(N__29409));
    Span4Mux_h I__5264 (
            .O(N__29409),
            .I(N__29405));
    InMux I__5263 (
            .O(N__29408),
            .I(N__29402));
    Odrv4 I__5262 (
            .O(N__29405),
            .I(\current_shift_inst.un38_control_input_0 ));
    LocalMux I__5261 (
            .O(N__29402),
            .I(\current_shift_inst.un38_control_input_0 ));
    InMux I__5260 (
            .O(N__29397),
            .I(N__29394));
    LocalMux I__5259 (
            .O(N__29394),
            .I(N__29391));
    Odrv4 I__5258 (
            .O(N__29391),
            .I(\current_shift_inst.un4_control_input_axb_2 ));
    InMux I__5257 (
            .O(N__29388),
            .I(N__29385));
    LocalMux I__5256 (
            .O(N__29385),
            .I(N__29381));
    InMux I__5255 (
            .O(N__29384),
            .I(N__29377));
    Span4Mux_h I__5254 (
            .O(N__29381),
            .I(N__29374));
    InMux I__5253 (
            .O(N__29380),
            .I(N__29371));
    LocalMux I__5252 (
            .O(N__29377),
            .I(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ));
    Odrv4 I__5251 (
            .O(N__29374),
            .I(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ));
    LocalMux I__5250 (
            .O(N__29371),
            .I(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ));
    InMux I__5249 (
            .O(N__29364),
            .I(\current_shift_inst.un4_control_input_cry_1 ));
    InMux I__5248 (
            .O(N__29361),
            .I(N__29358));
    LocalMux I__5247 (
            .O(N__29358),
            .I(N__29355));
    Odrv4 I__5246 (
            .O(N__29355),
            .I(\current_shift_inst.un4_control_input_axb_3 ));
    InMux I__5245 (
            .O(N__29352),
            .I(N__29349));
    LocalMux I__5244 (
            .O(N__29349),
            .I(N__29345));
    InMux I__5243 (
            .O(N__29348),
            .I(N__29341));
    Span4Mux_h I__5242 (
            .O(N__29345),
            .I(N__29338));
    InMux I__5241 (
            .O(N__29344),
            .I(N__29335));
    LocalMux I__5240 (
            .O(N__29341),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    Odrv4 I__5239 (
            .O(N__29338),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    LocalMux I__5238 (
            .O(N__29335),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    InMux I__5237 (
            .O(N__29328),
            .I(\current_shift_inst.un4_control_input_cry_2 ));
    InMux I__5236 (
            .O(N__29325),
            .I(N__29322));
    LocalMux I__5235 (
            .O(N__29322),
            .I(\current_shift_inst.un4_control_input_axb_4 ));
    InMux I__5234 (
            .O(N__29319),
            .I(N__29316));
    LocalMux I__5233 (
            .O(N__29316),
            .I(N__29313));
    Span4Mux_h I__5232 (
            .O(N__29313),
            .I(N__29309));
    InMux I__5231 (
            .O(N__29312),
            .I(N__29306));
    Odrv4 I__5230 (
            .O(N__29309),
            .I(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ));
    LocalMux I__5229 (
            .O(N__29306),
            .I(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ));
    InMux I__5228 (
            .O(N__29301),
            .I(\current_shift_inst.un4_control_input_cry_3 ));
    InMux I__5227 (
            .O(N__29298),
            .I(N__29295));
    LocalMux I__5226 (
            .O(N__29295),
            .I(\current_shift_inst.un4_control_input_axb_5 ));
    CascadeMux I__5225 (
            .O(N__29292),
            .I(N__29289));
    InMux I__5224 (
            .O(N__29289),
            .I(N__29286));
    LocalMux I__5223 (
            .O(N__29286),
            .I(N__29282));
    CascadeMux I__5222 (
            .O(N__29285),
            .I(N__29277));
    Span4Mux_v I__5221 (
            .O(N__29282),
            .I(N__29274));
    InMux I__5220 (
            .O(N__29281),
            .I(N__29269));
    InMux I__5219 (
            .O(N__29280),
            .I(N__29269));
    InMux I__5218 (
            .O(N__29277),
            .I(N__29266));
    Odrv4 I__5217 (
            .O(N__29274),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    LocalMux I__5216 (
            .O(N__29269),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    LocalMux I__5215 (
            .O(N__29266),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    InMux I__5214 (
            .O(N__29259),
            .I(\current_shift_inst.un4_control_input_cry_4 ));
    InMux I__5213 (
            .O(N__29256),
            .I(N__29253));
    LocalMux I__5212 (
            .O(N__29253),
            .I(\current_shift_inst.un4_control_input_axb_6 ));
    InMux I__5211 (
            .O(N__29250),
            .I(N__29245));
    InMux I__5210 (
            .O(N__29249),
            .I(N__29240));
    InMux I__5209 (
            .O(N__29248),
            .I(N__29240));
    LocalMux I__5208 (
            .O(N__29245),
            .I(N__29234));
    LocalMux I__5207 (
            .O(N__29240),
            .I(N__29234));
    InMux I__5206 (
            .O(N__29239),
            .I(N__29231));
    Odrv4 I__5205 (
            .O(N__29234),
            .I(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ));
    LocalMux I__5204 (
            .O(N__29231),
            .I(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ));
    InMux I__5203 (
            .O(N__29226),
            .I(\current_shift_inst.un4_control_input_cry_5 ));
    InMux I__5202 (
            .O(N__29223),
            .I(N__29220));
    LocalMux I__5201 (
            .O(N__29220),
            .I(\current_shift_inst.un4_control_input_axb_7 ));
    InMux I__5200 (
            .O(N__29217),
            .I(N__29211));
    InMux I__5199 (
            .O(N__29216),
            .I(N__29211));
    LocalMux I__5198 (
            .O(N__29211),
            .I(N__29207));
    InMux I__5197 (
            .O(N__29210),
            .I(N__29204));
    Span4Mux_h I__5196 (
            .O(N__29207),
            .I(N__29200));
    LocalMux I__5195 (
            .O(N__29204),
            .I(N__29197));
    InMux I__5194 (
            .O(N__29203),
            .I(N__29194));
    Odrv4 I__5193 (
            .O(N__29200),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    Odrv12 I__5192 (
            .O(N__29197),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    LocalMux I__5191 (
            .O(N__29194),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    InMux I__5190 (
            .O(N__29187),
            .I(\current_shift_inst.un4_control_input_cry_6 ));
    InMux I__5189 (
            .O(N__29184),
            .I(N__29181));
    LocalMux I__5188 (
            .O(N__29181),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ));
    InMux I__5187 (
            .O(N__29178),
            .I(N__29175));
    LocalMux I__5186 (
            .O(N__29175),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ));
    InMux I__5185 (
            .O(N__29172),
            .I(N__29168));
    InMux I__5184 (
            .O(N__29171),
            .I(N__29165));
    LocalMux I__5183 (
            .O(N__29168),
            .I(measured_delay_hc_27));
    LocalMux I__5182 (
            .O(N__29165),
            .I(measured_delay_hc_27));
    InMux I__5181 (
            .O(N__29160),
            .I(N__29157));
    LocalMux I__5180 (
            .O(N__29157),
            .I(N__29154));
    Odrv4 I__5179 (
            .O(N__29154),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4 ));
    CascadeMux I__5178 (
            .O(N__29151),
            .I(N__29148));
    InMux I__5177 (
            .O(N__29148),
            .I(N__29145));
    LocalMux I__5176 (
            .O(N__29145),
            .I(N__29142));
    Span4Mux_v I__5175 (
            .O(N__29142),
            .I(N__29139));
    Odrv4 I__5174 (
            .O(N__29139),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ));
    CascadeMux I__5173 (
            .O(N__29136),
            .I(N__29133));
    InMux I__5172 (
            .O(N__29133),
            .I(N__29126));
    InMux I__5171 (
            .O(N__29132),
            .I(N__29126));
    InMux I__5170 (
            .O(N__29131),
            .I(N__29123));
    LocalMux I__5169 (
            .O(N__29126),
            .I(N__29118));
    LocalMux I__5168 (
            .O(N__29123),
            .I(N__29118));
    Span4Mux_h I__5167 (
            .O(N__29118),
            .I(N__29114));
    InMux I__5166 (
            .O(N__29117),
            .I(N__29111));
    Odrv4 I__5165 (
            .O(N__29114),
            .I(\current_shift_inst.elapsed_time_ns_phase_6 ));
    LocalMux I__5164 (
            .O(N__29111),
            .I(\current_shift_inst.elapsed_time_ns_phase_6 ));
    CascadeMux I__5163 (
            .O(N__29106),
            .I(N__29103));
    InMux I__5162 (
            .O(N__29103),
            .I(N__29098));
    InMux I__5161 (
            .O(N__29102),
            .I(N__29093));
    InMux I__5160 (
            .O(N__29101),
            .I(N__29093));
    LocalMux I__5159 (
            .O(N__29098),
            .I(N__29088));
    LocalMux I__5158 (
            .O(N__29093),
            .I(N__29088));
    Span4Mux_h I__5157 (
            .O(N__29088),
            .I(N__29084));
    InMux I__5156 (
            .O(N__29087),
            .I(N__29081));
    Odrv4 I__5155 (
            .O(N__29084),
            .I(\current_shift_inst.elapsed_time_ns_phase_5 ));
    LocalMux I__5154 (
            .O(N__29081),
            .I(\current_shift_inst.elapsed_time_ns_phase_5 ));
    InMux I__5153 (
            .O(N__29076),
            .I(N__29073));
    LocalMux I__5152 (
            .O(N__29073),
            .I(N__29070));
    Odrv12 I__5151 (
            .O(N__29070),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ));
    InMux I__5150 (
            .O(N__29067),
            .I(N__29063));
    InMux I__5149 (
            .O(N__29066),
            .I(N__29060));
    LocalMux I__5148 (
            .O(N__29063),
            .I(measured_delay_hc_23));
    LocalMux I__5147 (
            .O(N__29060),
            .I(measured_delay_hc_23));
    CascadeMux I__5146 (
            .O(N__29055),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_3_cascade_ ));
    InMux I__5145 (
            .O(N__29052),
            .I(N__29046));
    InMux I__5144 (
            .O(N__29051),
            .I(N__29046));
    LocalMux I__5143 (
            .O(N__29046),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_14 ));
    InMux I__5142 (
            .O(N__29043),
            .I(N__29040));
    LocalMux I__5141 (
            .O(N__29040),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ));
    CascadeMux I__5140 (
            .O(N__29037),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt30_0_cascade_ ));
    InMux I__5139 (
            .O(N__29034),
            .I(N__29031));
    LocalMux I__5138 (
            .O(N__29031),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6 ));
    InMux I__5137 (
            .O(N__29028),
            .I(N__29025));
    LocalMux I__5136 (
            .O(N__29025),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_6 ));
    IoInMux I__5135 (
            .O(N__29022),
            .I(N__29019));
    LocalMux I__5134 (
            .O(N__29019),
            .I(N__29016));
    IoSpan4Mux I__5133 (
            .O(N__29016),
            .I(N__29013));
    IoSpan4Mux I__5132 (
            .O(N__29013),
            .I(N__29010));
    Span4Mux_s1_v I__5131 (
            .O(N__29010),
            .I(N__29007));
    Sp12to4 I__5130 (
            .O(N__29007),
            .I(N__29004));
    Span12Mux_s9_v I__5129 (
            .O(N__29004),
            .I(N__29001));
    Odrv12 I__5128 (
            .O(N__29001),
            .I(\current_shift_inst.timer_s1.N_187_i ));
    InMux I__5127 (
            .O(N__28998),
            .I(N__28995));
    LocalMux I__5126 (
            .O(N__28995),
            .I(N__28991));
    CascadeMux I__5125 (
            .O(N__28994),
            .I(N__28988));
    Span4Mux_v I__5124 (
            .O(N__28991),
            .I(N__28983));
    InMux I__5123 (
            .O(N__28988),
            .I(N__28977));
    InMux I__5122 (
            .O(N__28987),
            .I(N__28977));
    InMux I__5121 (
            .O(N__28986),
            .I(N__28974));
    Span4Mux_h I__5120 (
            .O(N__28983),
            .I(N__28971));
    InMux I__5119 (
            .O(N__28982),
            .I(N__28968));
    LocalMux I__5118 (
            .O(N__28977),
            .I(\current_shift_inst.phase_validZ0 ));
    LocalMux I__5117 (
            .O(N__28974),
            .I(\current_shift_inst.phase_validZ0 ));
    Odrv4 I__5116 (
            .O(N__28971),
            .I(\current_shift_inst.phase_validZ0 ));
    LocalMux I__5115 (
            .O(N__28968),
            .I(\current_shift_inst.phase_validZ0 ));
    CascadeMux I__5114 (
            .O(N__28959),
            .I(N__28955));
    InMux I__5113 (
            .O(N__28958),
            .I(N__28951));
    InMux I__5112 (
            .O(N__28955),
            .I(N__28948));
    InMux I__5111 (
            .O(N__28954),
            .I(N__28945));
    LocalMux I__5110 (
            .O(N__28951),
            .I(measured_delay_hc_20));
    LocalMux I__5109 (
            .O(N__28948),
            .I(measured_delay_hc_20));
    LocalMux I__5108 (
            .O(N__28945),
            .I(measured_delay_hc_20));
    InMux I__5107 (
            .O(N__28938),
            .I(N__28935));
    LocalMux I__5106 (
            .O(N__28935),
            .I(\current_shift_inst.z_5_27 ));
    InMux I__5105 (
            .O(N__28932),
            .I(N__28929));
    LocalMux I__5104 (
            .O(N__28929),
            .I(\current_shift_inst.z_5_28 ));
    CascadeMux I__5103 (
            .O(N__28926),
            .I(N__28923));
    InMux I__5102 (
            .O(N__28923),
            .I(N__28920));
    LocalMux I__5101 (
            .O(N__28920),
            .I(\current_shift_inst.z_5_29 ));
    CascadeMux I__5100 (
            .O(N__28917),
            .I(N__28914));
    InMux I__5099 (
            .O(N__28914),
            .I(N__28911));
    LocalMux I__5098 (
            .O(N__28911),
            .I(\current_shift_inst.z_5_30 ));
    InMux I__5097 (
            .O(N__28908),
            .I(N__28905));
    LocalMux I__5096 (
            .O(N__28905),
            .I(\current_shift_inst.z_5_cry_30_THRU_CO ));
    InMux I__5095 (
            .O(N__28902),
            .I(\current_shift_inst.z_cry_30 ));
    CascadeMux I__5094 (
            .O(N__28899),
            .I(N__28894));
    InMux I__5093 (
            .O(N__28898),
            .I(N__28889));
    InMux I__5092 (
            .O(N__28897),
            .I(N__28889));
    InMux I__5091 (
            .O(N__28894),
            .I(N__28886));
    LocalMux I__5090 (
            .O(N__28889),
            .I(N__28883));
    LocalMux I__5089 (
            .O(N__28886),
            .I(measured_delay_hc_21));
    Odrv4 I__5088 (
            .O(N__28883),
            .I(measured_delay_hc_21));
    CascadeMux I__5087 (
            .O(N__28878),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0_cascade_ ));
    InMux I__5086 (
            .O(N__28875),
            .I(N__28872));
    LocalMux I__5085 (
            .O(N__28872),
            .I(\current_shift_inst.z_5_19 ));
    CascadeMux I__5084 (
            .O(N__28869),
            .I(N__28866));
    InMux I__5083 (
            .O(N__28866),
            .I(N__28863));
    LocalMux I__5082 (
            .O(N__28863),
            .I(\current_shift_inst.z_5_20 ));
    InMux I__5081 (
            .O(N__28860),
            .I(N__28857));
    LocalMux I__5080 (
            .O(N__28857),
            .I(\current_shift_inst.z_5_21 ));
    InMux I__5079 (
            .O(N__28854),
            .I(N__28851));
    LocalMux I__5078 (
            .O(N__28851),
            .I(\current_shift_inst.z_5_22 ));
    InMux I__5077 (
            .O(N__28848),
            .I(N__28845));
    LocalMux I__5076 (
            .O(N__28845),
            .I(\current_shift_inst.z_5_23 ));
    InMux I__5075 (
            .O(N__28842),
            .I(N__28839));
    LocalMux I__5074 (
            .O(N__28839),
            .I(\current_shift_inst.z_5_24 ));
    CascadeMux I__5073 (
            .O(N__28836),
            .I(N__28833));
    InMux I__5072 (
            .O(N__28833),
            .I(N__28830));
    LocalMux I__5071 (
            .O(N__28830),
            .I(\current_shift_inst.z_5_25 ));
    InMux I__5070 (
            .O(N__28827),
            .I(N__28824));
    LocalMux I__5069 (
            .O(N__28824),
            .I(\current_shift_inst.z_5_26 ));
    InMux I__5068 (
            .O(N__28821),
            .I(N__28818));
    LocalMux I__5067 (
            .O(N__28818),
            .I(\current_shift_inst.z_5_10 ));
    InMux I__5066 (
            .O(N__28815),
            .I(N__28812));
    LocalMux I__5065 (
            .O(N__28812),
            .I(\current_shift_inst.z_5_11 ));
    InMux I__5064 (
            .O(N__28809),
            .I(N__28806));
    LocalMux I__5063 (
            .O(N__28806),
            .I(\current_shift_inst.z_5_12 ));
    InMux I__5062 (
            .O(N__28803),
            .I(N__28800));
    LocalMux I__5061 (
            .O(N__28800),
            .I(\current_shift_inst.z_5_13 ));
    InMux I__5060 (
            .O(N__28797),
            .I(N__28794));
    LocalMux I__5059 (
            .O(N__28794),
            .I(\current_shift_inst.z_5_14 ));
    InMux I__5058 (
            .O(N__28791),
            .I(N__28788));
    LocalMux I__5057 (
            .O(N__28788),
            .I(\current_shift_inst.z_5_15 ));
    InMux I__5056 (
            .O(N__28785),
            .I(N__28782));
    LocalMux I__5055 (
            .O(N__28782),
            .I(N__28779));
    Odrv4 I__5054 (
            .O(N__28779),
            .I(\current_shift_inst.z_5_16 ));
    InMux I__5053 (
            .O(N__28776),
            .I(N__28773));
    LocalMux I__5052 (
            .O(N__28773),
            .I(\current_shift_inst.z_5_17 ));
    InMux I__5051 (
            .O(N__28770),
            .I(N__28767));
    LocalMux I__5050 (
            .O(N__28767),
            .I(\current_shift_inst.z_5_18 ));
    CascadeMux I__5049 (
            .O(N__28764),
            .I(N__28761));
    InMux I__5048 (
            .O(N__28761),
            .I(N__28758));
    LocalMux I__5047 (
            .O(N__28758),
            .I(\current_shift_inst.z_5_2 ));
    CascadeMux I__5046 (
            .O(N__28755),
            .I(N__28752));
    InMux I__5045 (
            .O(N__28752),
            .I(N__28749));
    LocalMux I__5044 (
            .O(N__28749),
            .I(\current_shift_inst.z_5_3 ));
    InMux I__5043 (
            .O(N__28746),
            .I(N__28743));
    LocalMux I__5042 (
            .O(N__28743),
            .I(\current_shift_inst.z_5_4 ));
    CascadeMux I__5041 (
            .O(N__28740),
            .I(N__28737));
    InMux I__5040 (
            .O(N__28737),
            .I(N__28734));
    LocalMux I__5039 (
            .O(N__28734),
            .I(\current_shift_inst.z_5_5 ));
    CascadeMux I__5038 (
            .O(N__28731),
            .I(N__28728));
    InMux I__5037 (
            .O(N__28728),
            .I(N__28725));
    LocalMux I__5036 (
            .O(N__28725),
            .I(\current_shift_inst.z_5_6 ));
    InMux I__5035 (
            .O(N__28722),
            .I(N__28719));
    LocalMux I__5034 (
            .O(N__28719),
            .I(\current_shift_inst.z_5_7 ));
    InMux I__5033 (
            .O(N__28716),
            .I(N__28713));
    LocalMux I__5032 (
            .O(N__28713),
            .I(N__28710));
    Odrv4 I__5031 (
            .O(N__28710),
            .I(\current_shift_inst.z_5_8 ));
    InMux I__5030 (
            .O(N__28707),
            .I(N__28704));
    LocalMux I__5029 (
            .O(N__28704),
            .I(\current_shift_inst.z_5_9 ));
    InMux I__5028 (
            .O(N__28701),
            .I(N__28697));
    InMux I__5027 (
            .O(N__28700),
            .I(N__28694));
    LocalMux I__5026 (
            .O(N__28697),
            .I(N__28691));
    LocalMux I__5025 (
            .O(N__28694),
            .I(N__28688));
    Span4Mux_h I__5024 (
            .O(N__28691),
            .I(N__28684));
    Span4Mux_h I__5023 (
            .O(N__28688),
            .I(N__28681));
    InMux I__5022 (
            .O(N__28687),
            .I(N__28678));
    Odrv4 I__5021 (
            .O(N__28684),
            .I(\current_shift_inst.timer_phase.counterZ0Z_1 ));
    Odrv4 I__5020 (
            .O(N__28681),
            .I(\current_shift_inst.timer_phase.counterZ0Z_1 ));
    LocalMux I__5019 (
            .O(N__28678),
            .I(\current_shift_inst.timer_phase.counterZ0Z_1 ));
    InMux I__5018 (
            .O(N__28671),
            .I(N__28668));
    LocalMux I__5017 (
            .O(N__28668),
            .I(N__28665));
    Span4Mux_v I__5016 (
            .O(N__28665),
            .I(N__28662));
    Odrv4 I__5015 (
            .O(N__28662),
            .I(\current_shift_inst.N_1633_i ));
    InMux I__5014 (
            .O(N__28659),
            .I(N__28656));
    LocalMux I__5013 (
            .O(N__28656),
            .I(N__28652));
    InMux I__5012 (
            .O(N__28655),
            .I(N__28649));
    Span4Mux_h I__5011 (
            .O(N__28652),
            .I(N__28645));
    LocalMux I__5010 (
            .O(N__28649),
            .I(N__28642));
    InMux I__5009 (
            .O(N__28648),
            .I(N__28639));
    Odrv4 I__5008 (
            .O(N__28645),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    Odrv4 I__5007 (
            .O(N__28642),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    LocalMux I__5006 (
            .O(N__28639),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    CEMux I__5005 (
            .O(N__28632),
            .I(N__28617));
    CEMux I__5004 (
            .O(N__28631),
            .I(N__28617));
    CEMux I__5003 (
            .O(N__28630),
            .I(N__28617));
    CEMux I__5002 (
            .O(N__28629),
            .I(N__28617));
    CEMux I__5001 (
            .O(N__28628),
            .I(N__28617));
    GlobalMux I__5000 (
            .O(N__28617),
            .I(N__28614));
    gio2CtrlBuf I__4999 (
            .O(N__28614),
            .I(\current_shift_inst.timer_phase.N_188_i_g ));
    CascadeMux I__4998 (
            .O(N__28611),
            .I(N__28608));
    InMux I__4997 (
            .O(N__28608),
            .I(N__28605));
    LocalMux I__4996 (
            .O(N__28605),
            .I(N__28602));
    Span4Mux_v I__4995 (
            .O(N__28602),
            .I(N__28599));
    Odrv4 I__4994 (
            .O(N__28599),
            .I(\current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ));
    InMux I__4993 (
            .O(N__28596),
            .I(N__28590));
    InMux I__4992 (
            .O(N__28595),
            .I(N__28590));
    LocalMux I__4991 (
            .O(N__28590),
            .I(N__28586));
    CascadeMux I__4990 (
            .O(N__28589),
            .I(N__28583));
    Span4Mux_v I__4989 (
            .O(N__28586),
            .I(N__28580));
    InMux I__4988 (
            .O(N__28583),
            .I(N__28577));
    Odrv4 I__4987 (
            .O(N__28580),
            .I(\current_shift_inst.elapsed_time_ns_phase_3 ));
    LocalMux I__4986 (
            .O(N__28577),
            .I(\current_shift_inst.elapsed_time_ns_phase_3 ));
    CascadeMux I__4985 (
            .O(N__28572),
            .I(N__28567));
    InMux I__4984 (
            .O(N__28571),
            .I(N__28563));
    InMux I__4983 (
            .O(N__28570),
            .I(N__28560));
    InMux I__4982 (
            .O(N__28567),
            .I(N__28555));
    InMux I__4981 (
            .O(N__28566),
            .I(N__28555));
    LocalMux I__4980 (
            .O(N__28563),
            .I(N__28552));
    LocalMux I__4979 (
            .O(N__28560),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    LocalMux I__4978 (
            .O(N__28555),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    Odrv4 I__4977 (
            .O(N__28552),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    CascadeMux I__4976 (
            .O(N__28545),
            .I(N__28542));
    InMux I__4975 (
            .O(N__28542),
            .I(N__28539));
    LocalMux I__4974 (
            .O(N__28539),
            .I(N__28536));
    Span4Mux_v I__4973 (
            .O(N__28536),
            .I(N__28533));
    Odrv4 I__4972 (
            .O(N__28533),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ));
    CascadeMux I__4971 (
            .O(N__28530),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_ ));
    InMux I__4970 (
            .O(N__28527),
            .I(N__28524));
    LocalMux I__4969 (
            .O(N__28524),
            .I(N__28521));
    Span4Mux_h I__4968 (
            .O(N__28521),
            .I(N__28518));
    Odrv4 I__4967 (
            .O(N__28518),
            .I(\current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ));
    InMux I__4966 (
            .O(N__28515),
            .I(N__28511));
    CascadeMux I__4965 (
            .O(N__28514),
            .I(N__28508));
    LocalMux I__4964 (
            .O(N__28511),
            .I(N__28504));
    InMux I__4963 (
            .O(N__28508),
            .I(N__28499));
    InMux I__4962 (
            .O(N__28507),
            .I(N__28499));
    Span4Mux_h I__4961 (
            .O(N__28504),
            .I(N__28494));
    LocalMux I__4960 (
            .O(N__28499),
            .I(N__28494));
    Span4Mux_v I__4959 (
            .O(N__28494),
            .I(N__28490));
    InMux I__4958 (
            .O(N__28493),
            .I(N__28487));
    Odrv4 I__4957 (
            .O(N__28490),
            .I(\current_shift_inst.elapsed_time_ns_phase_4 ));
    LocalMux I__4956 (
            .O(N__28487),
            .I(\current_shift_inst.elapsed_time_ns_phase_4 ));
    CascadeMux I__4955 (
            .O(N__28482),
            .I(N__28479));
    InMux I__4954 (
            .O(N__28479),
            .I(N__28476));
    LocalMux I__4953 (
            .O(N__28476),
            .I(N__28473));
    Span4Mux_h I__4952 (
            .O(N__28473),
            .I(N__28470));
    Odrv4 I__4951 (
            .O(N__28470),
            .I(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ));
    CascadeMux I__4950 (
            .O(N__28467),
            .I(N__28464));
    InMux I__4949 (
            .O(N__28464),
            .I(N__28461));
    LocalMux I__4948 (
            .O(N__28461),
            .I(G_406));
    CascadeMux I__4947 (
            .O(N__28458),
            .I(N__28454));
    InMux I__4946 (
            .O(N__28457),
            .I(N__28447));
    InMux I__4945 (
            .O(N__28454),
            .I(N__28444));
    InMux I__4944 (
            .O(N__28453),
            .I(N__28435));
    InMux I__4943 (
            .O(N__28452),
            .I(N__28435));
    InMux I__4942 (
            .O(N__28451),
            .I(N__28435));
    InMux I__4941 (
            .O(N__28450),
            .I(N__28435));
    LocalMux I__4940 (
            .O(N__28447),
            .I(N__28430));
    LocalMux I__4939 (
            .O(N__28444),
            .I(N__28430));
    LocalMux I__4938 (
            .O(N__28435),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    Odrv4 I__4937 (
            .O(N__28430),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    CascadeMux I__4936 (
            .O(N__28425),
            .I(N__28422));
    InMux I__4935 (
            .O(N__28422),
            .I(N__28419));
    LocalMux I__4934 (
            .O(N__28419),
            .I(G_405));
    InMux I__4933 (
            .O(N__28416),
            .I(N__28409));
    InMux I__4932 (
            .O(N__28415),
            .I(N__28409));
    InMux I__4931 (
            .O(N__28414),
            .I(N__28406));
    LocalMux I__4930 (
            .O(N__28409),
            .I(N__28403));
    LocalMux I__4929 (
            .O(N__28406),
            .I(N__28400));
    Span4Mux_h I__4928 (
            .O(N__28403),
            .I(N__28394));
    Span4Mux_h I__4927 (
            .O(N__28400),
            .I(N__28394));
    InMux I__4926 (
            .O(N__28399),
            .I(N__28391));
    Odrv4 I__4925 (
            .O(N__28394),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    LocalMux I__4924 (
            .O(N__28391),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    CascadeMux I__4923 (
            .O(N__28386),
            .I(N__28383));
    InMux I__4922 (
            .O(N__28383),
            .I(N__28380));
    LocalMux I__4921 (
            .O(N__28380),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ));
    InMux I__4920 (
            .O(N__28377),
            .I(N__28368));
    InMux I__4919 (
            .O(N__28376),
            .I(N__28368));
    InMux I__4918 (
            .O(N__28375),
            .I(N__28368));
    LocalMux I__4917 (
            .O(N__28368),
            .I(N__28365));
    Span4Mux_h I__4916 (
            .O(N__28365),
            .I(N__28361));
    InMux I__4915 (
            .O(N__28364),
            .I(N__28358));
    Odrv4 I__4914 (
            .O(N__28361),
            .I(\current_shift_inst.elapsed_time_ns_phase_16 ));
    LocalMux I__4913 (
            .O(N__28358),
            .I(\current_shift_inst.elapsed_time_ns_phase_16 ));
    InMux I__4912 (
            .O(N__28353),
            .I(N__28350));
    LocalMux I__4911 (
            .O(N__28350),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ));
    InMux I__4910 (
            .O(N__28347),
            .I(N__28342));
    InMux I__4909 (
            .O(N__28346),
            .I(N__28339));
    InMux I__4908 (
            .O(N__28345),
            .I(N__28336));
    LocalMux I__4907 (
            .O(N__28342),
            .I(N__28331));
    LocalMux I__4906 (
            .O(N__28339),
            .I(N__28331));
    LocalMux I__4905 (
            .O(N__28336),
            .I(N__28325));
    Span4Mux_h I__4904 (
            .O(N__28331),
            .I(N__28325));
    InMux I__4903 (
            .O(N__28330),
            .I(N__28322));
    Span4Mux_v I__4902 (
            .O(N__28325),
            .I(N__28319));
    LocalMux I__4901 (
            .O(N__28322),
            .I(N__28316));
    Odrv4 I__4900 (
            .O(N__28319),
            .I(\current_shift_inst.elapsed_time_ns_phase_17 ));
    Odrv4 I__4899 (
            .O(N__28316),
            .I(\current_shift_inst.elapsed_time_ns_phase_17 ));
    CascadeMux I__4898 (
            .O(N__28311),
            .I(N__28308));
    InMux I__4897 (
            .O(N__28308),
            .I(N__28305));
    LocalMux I__4896 (
            .O(N__28305),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ));
    InMux I__4895 (
            .O(N__28302),
            .I(N__28297));
    InMux I__4894 (
            .O(N__28301),
            .I(N__28294));
    InMux I__4893 (
            .O(N__28300),
            .I(N__28291));
    LocalMux I__4892 (
            .O(N__28297),
            .I(N__28284));
    LocalMux I__4891 (
            .O(N__28294),
            .I(N__28284));
    LocalMux I__4890 (
            .O(N__28291),
            .I(N__28284));
    Span4Mux_v I__4889 (
            .O(N__28284),
            .I(N__28281));
    Span4Mux_v I__4888 (
            .O(N__28281),
            .I(N__28277));
    InMux I__4887 (
            .O(N__28280),
            .I(N__28274));
    Odrv4 I__4886 (
            .O(N__28277),
            .I(\current_shift_inst.elapsed_time_ns_phase_12 ));
    LocalMux I__4885 (
            .O(N__28274),
            .I(\current_shift_inst.elapsed_time_ns_phase_12 ));
    CascadeMux I__4884 (
            .O(N__28269),
            .I(N__28266));
    InMux I__4883 (
            .O(N__28266),
            .I(N__28263));
    LocalMux I__4882 (
            .O(N__28263),
            .I(N__28258));
    InMux I__4881 (
            .O(N__28262),
            .I(N__28253));
    InMux I__4880 (
            .O(N__28261),
            .I(N__28253));
    Span4Mux_h I__4879 (
            .O(N__28258),
            .I(N__28248));
    LocalMux I__4878 (
            .O(N__28253),
            .I(N__28248));
    Span4Mux_h I__4877 (
            .O(N__28248),
            .I(N__28244));
    InMux I__4876 (
            .O(N__28247),
            .I(N__28241));
    Odrv4 I__4875 (
            .O(N__28244),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    LocalMux I__4874 (
            .O(N__28241),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    InMux I__4873 (
            .O(N__28236),
            .I(N__28233));
    LocalMux I__4872 (
            .O(N__28233),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ));
    CascadeMux I__4871 (
            .O(N__28230),
            .I(N__28227));
    InMux I__4870 (
            .O(N__28227),
            .I(N__28224));
    LocalMux I__4869 (
            .O(N__28224),
            .I(N__28221));
    Span4Mux_v I__4868 (
            .O(N__28221),
            .I(N__28218));
    Odrv4 I__4867 (
            .O(N__28218),
            .I(\current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ));
    CascadeMux I__4866 (
            .O(N__28215),
            .I(N__28212));
    InMux I__4865 (
            .O(N__28212),
            .I(N__28209));
    LocalMux I__4864 (
            .O(N__28209),
            .I(N__28206));
    Odrv4 I__4863 (
            .O(N__28206),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ));
    InMux I__4862 (
            .O(N__28203),
            .I(N__28200));
    LocalMux I__4861 (
            .O(N__28200),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ));
    InMux I__4860 (
            .O(N__28197),
            .I(N__28188));
    InMux I__4859 (
            .O(N__28196),
            .I(N__28188));
    InMux I__4858 (
            .O(N__28195),
            .I(N__28188));
    LocalMux I__4857 (
            .O(N__28188),
            .I(N__28184));
    CascadeMux I__4856 (
            .O(N__28187),
            .I(N__28181));
    Span4Mux_h I__4855 (
            .O(N__28184),
            .I(N__28178));
    InMux I__4854 (
            .O(N__28181),
            .I(N__28175));
    Odrv4 I__4853 (
            .O(N__28178),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    LocalMux I__4852 (
            .O(N__28175),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    InMux I__4851 (
            .O(N__28170),
            .I(N__28167));
    LocalMux I__4850 (
            .O(N__28167),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ));
    CascadeMux I__4849 (
            .O(N__28164),
            .I(N__28161));
    InMux I__4848 (
            .O(N__28161),
            .I(N__28154));
    InMux I__4847 (
            .O(N__28160),
            .I(N__28154));
    InMux I__4846 (
            .O(N__28159),
            .I(N__28151));
    LocalMux I__4845 (
            .O(N__28154),
            .I(N__28148));
    LocalMux I__4844 (
            .O(N__28151),
            .I(N__28142));
    Span4Mux_h I__4843 (
            .O(N__28148),
            .I(N__28142));
    InMux I__4842 (
            .O(N__28147),
            .I(N__28139));
    Odrv4 I__4841 (
            .O(N__28142),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    LocalMux I__4840 (
            .O(N__28139),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    CascadeMux I__4839 (
            .O(N__28134),
            .I(N__28131));
    InMux I__4838 (
            .O(N__28131),
            .I(N__28128));
    LocalMux I__4837 (
            .O(N__28128),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ));
    InMux I__4836 (
            .O(N__28125),
            .I(N__28122));
    LocalMux I__4835 (
            .O(N__28122),
            .I(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ));
    InMux I__4834 (
            .O(N__28119),
            .I(N__28116));
    LocalMux I__4833 (
            .O(N__28116),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ));
    CascadeMux I__4832 (
            .O(N__28113),
            .I(N__28110));
    InMux I__4831 (
            .O(N__28110),
            .I(N__28107));
    LocalMux I__4830 (
            .O(N__28107),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI190J_15 ));
    CascadeMux I__4829 (
            .O(N__28104),
            .I(N__28101));
    InMux I__4828 (
            .O(N__28101),
            .I(N__28098));
    LocalMux I__4827 (
            .O(N__28098),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ));
    InMux I__4826 (
            .O(N__28095),
            .I(N__28086));
    InMux I__4825 (
            .O(N__28094),
            .I(N__28086));
    InMux I__4824 (
            .O(N__28093),
            .I(N__28086));
    LocalMux I__4823 (
            .O(N__28086),
            .I(N__28083));
    Span4Mux_h I__4822 (
            .O(N__28083),
            .I(N__28079));
    InMux I__4821 (
            .O(N__28082),
            .I(N__28076));
    Odrv4 I__4820 (
            .O(N__28079),
            .I(\current_shift_inst.elapsed_time_ns_phase_15 ));
    LocalMux I__4819 (
            .O(N__28076),
            .I(\current_shift_inst.elapsed_time_ns_phase_15 ));
    InMux I__4818 (
            .O(N__28071),
            .I(N__28068));
    LocalMux I__4817 (
            .O(N__28068),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ));
    CascadeMux I__4816 (
            .O(N__28065),
            .I(N__28062));
    InMux I__4815 (
            .O(N__28062),
            .I(N__28059));
    LocalMux I__4814 (
            .O(N__28059),
            .I(N__28056));
    Odrv4 I__4813 (
            .O(N__28056),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ));
    CascadeMux I__4812 (
            .O(N__28053),
            .I(N__28050));
    InMux I__4811 (
            .O(N__28050),
            .I(N__28043));
    InMux I__4810 (
            .O(N__28049),
            .I(N__28043));
    InMux I__4809 (
            .O(N__28048),
            .I(N__28040));
    LocalMux I__4808 (
            .O(N__28043),
            .I(N__28037));
    LocalMux I__4807 (
            .O(N__28040),
            .I(N__28032));
    Span4Mux_h I__4806 (
            .O(N__28037),
            .I(N__28032));
    Sp12to4 I__4805 (
            .O(N__28032),
            .I(N__28028));
    InMux I__4804 (
            .O(N__28031),
            .I(N__28025));
    Odrv12 I__4803 (
            .O(N__28028),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    LocalMux I__4802 (
            .O(N__28025),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    InMux I__4801 (
            .O(N__28020),
            .I(N__28017));
    LocalMux I__4800 (
            .O(N__28017),
            .I(N__28014));
    Odrv4 I__4799 (
            .O(N__28014),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ));
    InMux I__4798 (
            .O(N__28011),
            .I(N__28008));
    LocalMux I__4797 (
            .O(N__28008),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ));
    CascadeMux I__4796 (
            .O(N__28005),
            .I(N__28002));
    InMux I__4795 (
            .O(N__28002),
            .I(N__27999));
    LocalMux I__4794 (
            .O(N__27999),
            .I(N__27996));
    Odrv4 I__4793 (
            .O(N__27996),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ));
    CascadeMux I__4792 (
            .O(N__27993),
            .I(N__27990));
    InMux I__4791 (
            .O(N__27990),
            .I(N__27987));
    LocalMux I__4790 (
            .O(N__27987),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ));
    CascadeMux I__4789 (
            .O(N__27984),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_5_cascade_ ));
    CascadeMux I__4788 (
            .O(N__27981),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_ ));
    InMux I__4787 (
            .O(N__27978),
            .I(N__27975));
    LocalMux I__4786 (
            .O(N__27975),
            .I(N__27972));
    Odrv4 I__4785 (
            .O(N__27972),
            .I(il_min_comp1_D1));
    CascadeMux I__4784 (
            .O(N__27969),
            .I(N__27966));
    InMux I__4783 (
            .O(N__27966),
            .I(N__27961));
    InMux I__4782 (
            .O(N__27965),
            .I(N__27956));
    InMux I__4781 (
            .O(N__27964),
            .I(N__27956));
    LocalMux I__4780 (
            .O(N__27961),
            .I(measured_delay_hc_22));
    LocalMux I__4779 (
            .O(N__27956),
            .I(measured_delay_hc_22));
    CascadeMux I__4778 (
            .O(N__27951),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_ ));
    InMux I__4777 (
            .O(N__27948),
            .I(\current_shift_inst.z_5_cry_25 ));
    CascadeMux I__4776 (
            .O(N__27945),
            .I(N__27941));
    InMux I__4775 (
            .O(N__27944),
            .I(N__27933));
    InMux I__4774 (
            .O(N__27941),
            .I(N__27933));
    InMux I__4773 (
            .O(N__27940),
            .I(N__27933));
    LocalMux I__4772 (
            .O(N__27933),
            .I(N__27930));
    Span4Mux_h I__4771 (
            .O(N__27930),
            .I(N__27926));
    InMux I__4770 (
            .O(N__27929),
            .I(N__27923));
    Odrv4 I__4769 (
            .O(N__27926),
            .I(\current_shift_inst.elapsed_time_ns_phase_27 ));
    LocalMux I__4768 (
            .O(N__27923),
            .I(\current_shift_inst.elapsed_time_ns_phase_27 ));
    InMux I__4767 (
            .O(N__27918),
            .I(\current_shift_inst.z_5_cry_26 ));
    InMux I__4766 (
            .O(N__27915),
            .I(N__27906));
    InMux I__4765 (
            .O(N__27914),
            .I(N__27906));
    InMux I__4764 (
            .O(N__27913),
            .I(N__27906));
    LocalMux I__4763 (
            .O(N__27906),
            .I(N__27903));
    Span4Mux_h I__4762 (
            .O(N__27903),
            .I(N__27899));
    InMux I__4761 (
            .O(N__27902),
            .I(N__27896));
    Odrv4 I__4760 (
            .O(N__27899),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    LocalMux I__4759 (
            .O(N__27896),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    InMux I__4758 (
            .O(N__27891),
            .I(\current_shift_inst.z_5_cry_27 ));
    CascadeMux I__4757 (
            .O(N__27888),
            .I(N__27884));
    InMux I__4756 (
            .O(N__27887),
            .I(N__27879));
    InMux I__4755 (
            .O(N__27884),
            .I(N__27879));
    LocalMux I__4754 (
            .O(N__27879),
            .I(N__27876));
    Span4Mux_h I__4753 (
            .O(N__27876),
            .I(N__27872));
    InMux I__4752 (
            .O(N__27875),
            .I(N__27869));
    Odrv4 I__4751 (
            .O(N__27872),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    LocalMux I__4750 (
            .O(N__27869),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    InMux I__4749 (
            .O(N__27864),
            .I(\current_shift_inst.z_5_cry_28 ));
    CascadeMux I__4748 (
            .O(N__27861),
            .I(N__27854));
    CascadeMux I__4747 (
            .O(N__27860),
            .I(N__27851));
    CascadeMux I__4746 (
            .O(N__27859),
            .I(N__27848));
    CascadeMux I__4745 (
            .O(N__27858),
            .I(N__27845));
    CascadeMux I__4744 (
            .O(N__27857),
            .I(N__27842));
    InMux I__4743 (
            .O(N__27854),
            .I(N__27823));
    InMux I__4742 (
            .O(N__27851),
            .I(N__27814));
    InMux I__4741 (
            .O(N__27848),
            .I(N__27814));
    InMux I__4740 (
            .O(N__27845),
            .I(N__27814));
    InMux I__4739 (
            .O(N__27842),
            .I(N__27814));
    CascadeMux I__4738 (
            .O(N__27841),
            .I(N__27811));
    CascadeMux I__4737 (
            .O(N__27840),
            .I(N__27808));
    CascadeMux I__4736 (
            .O(N__27839),
            .I(N__27805));
    CascadeMux I__4735 (
            .O(N__27838),
            .I(N__27802));
    InMux I__4734 (
            .O(N__27837),
            .I(N__27791));
    InMux I__4733 (
            .O(N__27836),
            .I(N__27791));
    InMux I__4732 (
            .O(N__27835),
            .I(N__27791));
    InMux I__4731 (
            .O(N__27834),
            .I(N__27788));
    InMux I__4730 (
            .O(N__27833),
            .I(N__27779));
    InMux I__4729 (
            .O(N__27832),
            .I(N__27779));
    InMux I__4728 (
            .O(N__27831),
            .I(N__27779));
    InMux I__4727 (
            .O(N__27830),
            .I(N__27779));
    CascadeMux I__4726 (
            .O(N__27829),
            .I(N__27769));
    CascadeMux I__4725 (
            .O(N__27828),
            .I(N__27766));
    CascadeMux I__4724 (
            .O(N__27827),
            .I(N__27763));
    CascadeMux I__4723 (
            .O(N__27826),
            .I(N__27760));
    LocalMux I__4722 (
            .O(N__27823),
            .I(N__27755));
    LocalMux I__4721 (
            .O(N__27814),
            .I(N__27755));
    InMux I__4720 (
            .O(N__27811),
            .I(N__27746));
    InMux I__4719 (
            .O(N__27808),
            .I(N__27746));
    InMux I__4718 (
            .O(N__27805),
            .I(N__27746));
    InMux I__4717 (
            .O(N__27802),
            .I(N__27746));
    CascadeMux I__4716 (
            .O(N__27801),
            .I(N__27743));
    CascadeMux I__4715 (
            .O(N__27800),
            .I(N__27740));
    CascadeMux I__4714 (
            .O(N__27799),
            .I(N__27737));
    CascadeMux I__4713 (
            .O(N__27798),
            .I(N__27734));
    LocalMux I__4712 (
            .O(N__27791),
            .I(N__27731));
    LocalMux I__4711 (
            .O(N__27788),
            .I(N__27726));
    LocalMux I__4710 (
            .O(N__27779),
            .I(N__27726));
    InMux I__4709 (
            .O(N__27778),
            .I(N__27723));
    CascadeMux I__4708 (
            .O(N__27777),
            .I(N__27720));
    CascadeMux I__4707 (
            .O(N__27776),
            .I(N__27717));
    CascadeMux I__4706 (
            .O(N__27775),
            .I(N__27706));
    CascadeMux I__4705 (
            .O(N__27774),
            .I(N__27702));
    CascadeMux I__4704 (
            .O(N__27773),
            .I(N__27699));
    CascadeMux I__4703 (
            .O(N__27772),
            .I(N__27695));
    InMux I__4702 (
            .O(N__27769),
            .I(N__27686));
    InMux I__4701 (
            .O(N__27766),
            .I(N__27686));
    InMux I__4700 (
            .O(N__27763),
            .I(N__27686));
    InMux I__4699 (
            .O(N__27760),
            .I(N__27686));
    Span4Mux_v I__4698 (
            .O(N__27755),
            .I(N__27681));
    LocalMux I__4697 (
            .O(N__27746),
            .I(N__27681));
    InMux I__4696 (
            .O(N__27743),
            .I(N__27672));
    InMux I__4695 (
            .O(N__27740),
            .I(N__27672));
    InMux I__4694 (
            .O(N__27737),
            .I(N__27672));
    InMux I__4693 (
            .O(N__27734),
            .I(N__27672));
    Span4Mux_v I__4692 (
            .O(N__27731),
            .I(N__27659));
    Span4Mux_v I__4691 (
            .O(N__27726),
            .I(N__27659));
    LocalMux I__4690 (
            .O(N__27723),
            .I(N__27659));
    InMux I__4689 (
            .O(N__27720),
            .I(N__27656));
    InMux I__4688 (
            .O(N__27717),
            .I(N__27651));
    InMux I__4687 (
            .O(N__27716),
            .I(N__27651));
    InMux I__4686 (
            .O(N__27715),
            .I(N__27644));
    InMux I__4685 (
            .O(N__27714),
            .I(N__27644));
    InMux I__4684 (
            .O(N__27713),
            .I(N__27644));
    InMux I__4683 (
            .O(N__27712),
            .I(N__27635));
    InMux I__4682 (
            .O(N__27711),
            .I(N__27635));
    InMux I__4681 (
            .O(N__27710),
            .I(N__27635));
    InMux I__4680 (
            .O(N__27709),
            .I(N__27635));
    InMux I__4679 (
            .O(N__27706),
            .I(N__27622));
    InMux I__4678 (
            .O(N__27705),
            .I(N__27622));
    InMux I__4677 (
            .O(N__27702),
            .I(N__27622));
    InMux I__4676 (
            .O(N__27699),
            .I(N__27622));
    InMux I__4675 (
            .O(N__27698),
            .I(N__27622));
    InMux I__4674 (
            .O(N__27695),
            .I(N__27622));
    LocalMux I__4673 (
            .O(N__27686),
            .I(N__27619));
    Span4Mux_h I__4672 (
            .O(N__27681),
            .I(N__27614));
    LocalMux I__4671 (
            .O(N__27672),
            .I(N__27614));
    CascadeMux I__4670 (
            .O(N__27671),
            .I(N__27611));
    CascadeMux I__4669 (
            .O(N__27670),
            .I(N__27608));
    CascadeMux I__4668 (
            .O(N__27669),
            .I(N__27605));
    CascadeMux I__4667 (
            .O(N__27668),
            .I(N__27602));
    CascadeMux I__4666 (
            .O(N__27667),
            .I(N__27599));
    CascadeMux I__4665 (
            .O(N__27666),
            .I(N__27596));
    Span4Mux_v I__4664 (
            .O(N__27659),
            .I(N__27592));
    LocalMux I__4663 (
            .O(N__27656),
            .I(N__27587));
    LocalMux I__4662 (
            .O(N__27651),
            .I(N__27587));
    LocalMux I__4661 (
            .O(N__27644),
            .I(N__27582));
    LocalMux I__4660 (
            .O(N__27635),
            .I(N__27582));
    LocalMux I__4659 (
            .O(N__27622),
            .I(N__27579));
    Span4Mux_v I__4658 (
            .O(N__27619),
            .I(N__27574));
    Span4Mux_v I__4657 (
            .O(N__27614),
            .I(N__27574));
    InMux I__4656 (
            .O(N__27611),
            .I(N__27567));
    InMux I__4655 (
            .O(N__27608),
            .I(N__27567));
    InMux I__4654 (
            .O(N__27605),
            .I(N__27567));
    InMux I__4653 (
            .O(N__27602),
            .I(N__27560));
    InMux I__4652 (
            .O(N__27599),
            .I(N__27560));
    InMux I__4651 (
            .O(N__27596),
            .I(N__27560));
    InMux I__4650 (
            .O(N__27595),
            .I(N__27557));
    Sp12to4 I__4649 (
            .O(N__27592),
            .I(N__27553));
    Span4Mux_v I__4648 (
            .O(N__27587),
            .I(N__27548));
    Span4Mux_s2_h I__4647 (
            .O(N__27582),
            .I(N__27548));
    Span4Mux_v I__4646 (
            .O(N__27579),
            .I(N__27539));
    Span4Mux_v I__4645 (
            .O(N__27574),
            .I(N__27539));
    LocalMux I__4644 (
            .O(N__27567),
            .I(N__27539));
    LocalMux I__4643 (
            .O(N__27560),
            .I(N__27539));
    LocalMux I__4642 (
            .O(N__27557),
            .I(N__27536));
    InMux I__4641 (
            .O(N__27556),
            .I(N__27532));
    Span12Mux_h I__4640 (
            .O(N__27553),
            .I(N__27526));
    Sp12to4 I__4639 (
            .O(N__27548),
            .I(N__27526));
    Sp12to4 I__4638 (
            .O(N__27539),
            .I(N__27523));
    Span12Mux_s3_h I__4637 (
            .O(N__27536),
            .I(N__27520));
    InMux I__4636 (
            .O(N__27535),
            .I(N__27517));
    LocalMux I__4635 (
            .O(N__27532),
            .I(N__27514));
    InMux I__4634 (
            .O(N__27531),
            .I(N__27511));
    Span12Mux_v I__4633 (
            .O(N__27526),
            .I(N__27508));
    Span12Mux_v I__4632 (
            .O(N__27523),
            .I(N__27501));
    Span12Mux_h I__4631 (
            .O(N__27520),
            .I(N__27501));
    LocalMux I__4630 (
            .O(N__27517),
            .I(N__27501));
    Span4Mux_s1_v I__4629 (
            .O(N__27514),
            .I(N__27496));
    LocalMux I__4628 (
            .O(N__27511),
            .I(N__27496));
    Odrv12 I__4627 (
            .O(N__27508),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4626 (
            .O(N__27501),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4625 (
            .O(N__27496),
            .I(CONSTANT_ONE_NET));
    InMux I__4624 (
            .O(N__27489),
            .I(\current_shift_inst.z_5_cry_29 ));
    InMux I__4623 (
            .O(N__27486),
            .I(\current_shift_inst.z_5_cry_30 ));
    InMux I__4622 (
            .O(N__27483),
            .I(N__27480));
    LocalMux I__4621 (
            .O(N__27480),
            .I(N__27477));
    Span4Mux_h I__4620 (
            .O(N__27477),
            .I(N__27474));
    Odrv4 I__4619 (
            .O(N__27474),
            .I(il_min_comp2_D1));
    InMux I__4618 (
            .O(N__27471),
            .I(N__27468));
    LocalMux I__4617 (
            .O(N__27468),
            .I(N__27462));
    InMux I__4616 (
            .O(N__27467),
            .I(N__27457));
    InMux I__4615 (
            .O(N__27466),
            .I(N__27457));
    InMux I__4614 (
            .O(N__27465),
            .I(N__27454));
    Span4Mux_h I__4613 (
            .O(N__27462),
            .I(N__27449));
    LocalMux I__4612 (
            .O(N__27457),
            .I(N__27449));
    LocalMux I__4611 (
            .O(N__27454),
            .I(N__27446));
    Odrv4 I__4610 (
            .O(N__27449),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    Odrv4 I__4609 (
            .O(N__27446),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    InMux I__4608 (
            .O(N__27441),
            .I(\current_shift_inst.z_5_cry_17 ));
    CascadeMux I__4607 (
            .O(N__27438),
            .I(N__27434));
    InMux I__4606 (
            .O(N__27437),
            .I(N__27426));
    InMux I__4605 (
            .O(N__27434),
            .I(N__27426));
    InMux I__4604 (
            .O(N__27433),
            .I(N__27426));
    LocalMux I__4603 (
            .O(N__27426),
            .I(N__27423));
    Span4Mux_h I__4602 (
            .O(N__27423),
            .I(N__27419));
    InMux I__4601 (
            .O(N__27422),
            .I(N__27416));
    Odrv4 I__4600 (
            .O(N__27419),
            .I(\current_shift_inst.elapsed_time_ns_phase_19 ));
    LocalMux I__4599 (
            .O(N__27416),
            .I(\current_shift_inst.elapsed_time_ns_phase_19 ));
    InMux I__4598 (
            .O(N__27411),
            .I(\current_shift_inst.z_5_cry_18 ));
    InMux I__4597 (
            .O(N__27408),
            .I(N__27399));
    InMux I__4596 (
            .O(N__27407),
            .I(N__27399));
    InMux I__4595 (
            .O(N__27406),
            .I(N__27399));
    LocalMux I__4594 (
            .O(N__27399),
            .I(N__27396));
    Span4Mux_h I__4593 (
            .O(N__27396),
            .I(N__27392));
    InMux I__4592 (
            .O(N__27395),
            .I(N__27389));
    Odrv4 I__4591 (
            .O(N__27392),
            .I(\current_shift_inst.elapsed_time_ns_phase_20 ));
    LocalMux I__4590 (
            .O(N__27389),
            .I(\current_shift_inst.elapsed_time_ns_phase_20 ));
    InMux I__4589 (
            .O(N__27384),
            .I(\current_shift_inst.z_5_cry_19 ));
    CascadeMux I__4588 (
            .O(N__27381),
            .I(N__27376));
    InMux I__4587 (
            .O(N__27380),
            .I(N__27373));
    InMux I__4586 (
            .O(N__27379),
            .I(N__27368));
    InMux I__4585 (
            .O(N__27376),
            .I(N__27368));
    LocalMux I__4584 (
            .O(N__27373),
            .I(N__27363));
    LocalMux I__4583 (
            .O(N__27368),
            .I(N__27363));
    Span4Mux_h I__4582 (
            .O(N__27363),
            .I(N__27359));
    InMux I__4581 (
            .O(N__27362),
            .I(N__27356));
    Odrv4 I__4580 (
            .O(N__27359),
            .I(\current_shift_inst.elapsed_time_ns_phase_21 ));
    LocalMux I__4579 (
            .O(N__27356),
            .I(\current_shift_inst.elapsed_time_ns_phase_21 ));
    InMux I__4578 (
            .O(N__27351),
            .I(\current_shift_inst.z_5_cry_20 ));
    InMux I__4577 (
            .O(N__27348),
            .I(\current_shift_inst.z_5_cry_21 ));
    InMux I__4576 (
            .O(N__27345),
            .I(\current_shift_inst.z_5_cry_22 ));
    InMux I__4575 (
            .O(N__27342),
            .I(\current_shift_inst.z_5_cry_23 ));
    InMux I__4574 (
            .O(N__27339),
            .I(bfn_9_21_0_));
    InMux I__4573 (
            .O(N__27336),
            .I(N__27327));
    InMux I__4572 (
            .O(N__27335),
            .I(N__27327));
    InMux I__4571 (
            .O(N__27334),
            .I(N__27327));
    LocalMux I__4570 (
            .O(N__27327),
            .I(N__27323));
    InMux I__4569 (
            .O(N__27326),
            .I(N__27320));
    Span4Mux_h I__4568 (
            .O(N__27323),
            .I(N__27317));
    LocalMux I__4567 (
            .O(N__27320),
            .I(N__27314));
    Odrv4 I__4566 (
            .O(N__27317),
            .I(\current_shift_inst.elapsed_time_ns_phase_9 ));
    Odrv4 I__4565 (
            .O(N__27314),
            .I(\current_shift_inst.elapsed_time_ns_phase_9 ));
    InMux I__4564 (
            .O(N__27309),
            .I(bfn_9_19_0_));
    InMux I__4563 (
            .O(N__27306),
            .I(N__27297));
    InMux I__4562 (
            .O(N__27305),
            .I(N__27297));
    InMux I__4561 (
            .O(N__27304),
            .I(N__27297));
    LocalMux I__4560 (
            .O(N__27297),
            .I(N__27293));
    InMux I__4559 (
            .O(N__27296),
            .I(N__27290));
    Span4Mux_h I__4558 (
            .O(N__27293),
            .I(N__27287));
    LocalMux I__4557 (
            .O(N__27290),
            .I(N__27284));
    Odrv4 I__4556 (
            .O(N__27287),
            .I(\current_shift_inst.elapsed_time_ns_phase_10 ));
    Odrv4 I__4555 (
            .O(N__27284),
            .I(\current_shift_inst.elapsed_time_ns_phase_10 ));
    InMux I__4554 (
            .O(N__27279),
            .I(\current_shift_inst.z_5_cry_9 ));
    InMux I__4553 (
            .O(N__27276),
            .I(\current_shift_inst.z_5_cry_10 ));
    InMux I__4552 (
            .O(N__27273),
            .I(\current_shift_inst.z_5_cry_11 ));
    InMux I__4551 (
            .O(N__27270),
            .I(\current_shift_inst.z_5_cry_12 ));
    InMux I__4550 (
            .O(N__27267),
            .I(\current_shift_inst.z_5_cry_13 ));
    InMux I__4549 (
            .O(N__27264),
            .I(\current_shift_inst.z_5_cry_14 ));
    InMux I__4548 (
            .O(N__27261),
            .I(\current_shift_inst.z_5_cry_15 ));
    InMux I__4547 (
            .O(N__27258),
            .I(bfn_9_20_0_));
    CascadeMux I__4546 (
            .O(N__27255),
            .I(N__27252));
    InMux I__4545 (
            .O(N__27252),
            .I(N__27249));
    LocalMux I__4544 (
            .O(N__27249),
            .I(\current_shift_inst.control_input_1_cry_24_THRU_CO ));
    InMux I__4543 (
            .O(N__27246),
            .I(bfn_9_17_0_));
    CascadeMux I__4542 (
            .O(N__27243),
            .I(N__27240));
    InMux I__4541 (
            .O(N__27240),
            .I(N__27234));
    CascadeMux I__4540 (
            .O(N__27239),
            .I(N__27229));
    CascadeMux I__4539 (
            .O(N__27238),
            .I(N__27226));
    CascadeMux I__4538 (
            .O(N__27237),
            .I(N__27222));
    LocalMux I__4537 (
            .O(N__27234),
            .I(N__27218));
    InMux I__4536 (
            .O(N__27233),
            .I(N__27215));
    InMux I__4535 (
            .O(N__27232),
            .I(N__27202));
    InMux I__4534 (
            .O(N__27229),
            .I(N__27202));
    InMux I__4533 (
            .O(N__27226),
            .I(N__27202));
    InMux I__4532 (
            .O(N__27225),
            .I(N__27202));
    InMux I__4531 (
            .O(N__27222),
            .I(N__27202));
    InMux I__4530 (
            .O(N__27221),
            .I(N__27202));
    Span4Mux_h I__4529 (
            .O(N__27218),
            .I(N__27199));
    LocalMux I__4528 (
            .O(N__27215),
            .I(N__27194));
    LocalMux I__4527 (
            .O(N__27202),
            .I(N__27194));
    Span4Mux_h I__4526 (
            .O(N__27199),
            .I(N__27189));
    Span4Mux_h I__4525 (
            .O(N__27194),
            .I(N__27189));
    Odrv4 I__4524 (
            .O(N__27189),
            .I(\current_shift_inst.control_inputZ0Z_25 ));
    CEMux I__4523 (
            .O(N__27186),
            .I(N__27181));
    CEMux I__4522 (
            .O(N__27185),
            .I(N__27178));
    CEMux I__4521 (
            .O(N__27184),
            .I(N__27175));
    LocalMux I__4520 (
            .O(N__27181),
            .I(N__27171));
    LocalMux I__4519 (
            .O(N__27178),
            .I(N__27166));
    LocalMux I__4518 (
            .O(N__27175),
            .I(N__27166));
    CEMux I__4517 (
            .O(N__27174),
            .I(N__27163));
    Span4Mux_v I__4516 (
            .O(N__27171),
            .I(N__27155));
    Span4Mux_v I__4515 (
            .O(N__27166),
            .I(N__27155));
    LocalMux I__4514 (
            .O(N__27163),
            .I(N__27155));
    CEMux I__4513 (
            .O(N__27162),
            .I(N__27152));
    Span4Mux_v I__4512 (
            .O(N__27155),
            .I(N__27149));
    LocalMux I__4511 (
            .O(N__27152),
            .I(N__27146));
    Span4Mux_v I__4510 (
            .O(N__27149),
            .I(N__27143));
    Span4Mux_v I__4509 (
            .O(N__27146),
            .I(N__27140));
    Odrv4 I__4508 (
            .O(N__27143),
            .I(\current_shift_inst.phase_valid_RNISLORZ0Z2 ));
    Odrv4 I__4507 (
            .O(N__27140),
            .I(\current_shift_inst.phase_valid_RNISLORZ0Z2 ));
    InMux I__4506 (
            .O(N__27135),
            .I(\current_shift_inst.z_5_cry_1 ));
    InMux I__4505 (
            .O(N__27132),
            .I(\current_shift_inst.z_5_cry_2 ));
    InMux I__4504 (
            .O(N__27129),
            .I(\current_shift_inst.z_5_cry_3 ));
    InMux I__4503 (
            .O(N__27126),
            .I(\current_shift_inst.z_5_cry_4 ));
    InMux I__4502 (
            .O(N__27123),
            .I(\current_shift_inst.z_5_cry_5 ));
    InMux I__4501 (
            .O(N__27120),
            .I(\current_shift_inst.z_5_cry_6 ));
    InMux I__4500 (
            .O(N__27117),
            .I(\current_shift_inst.z_5_cry_7 ));
    CascadeMux I__4499 (
            .O(N__27114),
            .I(N__27111));
    InMux I__4498 (
            .O(N__27111),
            .I(N__27108));
    LocalMux I__4497 (
            .O(N__27108),
            .I(N__27105));
    Span4Mux_h I__4496 (
            .O(N__27105),
            .I(N__27102));
    Odrv4 I__4495 (
            .O(N__27102),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ));
    InMux I__4494 (
            .O(N__27099),
            .I(N__27096));
    LocalMux I__4493 (
            .O(N__27096),
            .I(\current_shift_inst.control_input_1_axb_17 ));
    InMux I__4492 (
            .O(N__27093),
            .I(bfn_9_16_0_));
    InMux I__4491 (
            .O(N__27090),
            .I(N__27087));
    LocalMux I__4490 (
            .O(N__27087),
            .I(\current_shift_inst.control_input_1_axb_18 ));
    InMux I__4489 (
            .O(N__27084),
            .I(\current_shift_inst.un38_control_input_0_cry_23 ));
    InMux I__4488 (
            .O(N__27081),
            .I(N__27078));
    LocalMux I__4487 (
            .O(N__27078),
            .I(\current_shift_inst.control_input_1_axb_19 ));
    InMux I__4486 (
            .O(N__27075),
            .I(\current_shift_inst.un38_control_input_0_cry_24 ));
    InMux I__4485 (
            .O(N__27072),
            .I(N__27069));
    LocalMux I__4484 (
            .O(N__27069),
            .I(\current_shift_inst.control_input_1_axb_20 ));
    InMux I__4483 (
            .O(N__27066),
            .I(\current_shift_inst.un38_control_input_0_cry_25 ));
    InMux I__4482 (
            .O(N__27063),
            .I(N__27060));
    LocalMux I__4481 (
            .O(N__27060),
            .I(N__27057));
    Odrv4 I__4480 (
            .O(N__27057),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ));
    InMux I__4479 (
            .O(N__27054),
            .I(N__27051));
    LocalMux I__4478 (
            .O(N__27051),
            .I(\current_shift_inst.control_input_1_axb_21 ));
    InMux I__4477 (
            .O(N__27048),
            .I(\current_shift_inst.un38_control_input_0_cry_26 ));
    InMux I__4476 (
            .O(N__27045),
            .I(N__27042));
    LocalMux I__4475 (
            .O(N__27042),
            .I(N__27039));
    Odrv4 I__4474 (
            .O(N__27039),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ));
    CascadeMux I__4473 (
            .O(N__27036),
            .I(N__27033));
    InMux I__4472 (
            .O(N__27033),
            .I(N__27030));
    LocalMux I__4471 (
            .O(N__27030),
            .I(N__27027));
    Odrv4 I__4470 (
            .O(N__27027),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ));
    InMux I__4469 (
            .O(N__27024),
            .I(N__27021));
    LocalMux I__4468 (
            .O(N__27021),
            .I(\current_shift_inst.control_input_1_axb_22 ));
    InMux I__4467 (
            .O(N__27018),
            .I(\current_shift_inst.un38_control_input_0_cry_27 ));
    InMux I__4466 (
            .O(N__27015),
            .I(N__27012));
    LocalMux I__4465 (
            .O(N__27012),
            .I(N__27009));
    Odrv12 I__4464 (
            .O(N__27009),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ));
    CascadeMux I__4463 (
            .O(N__27006),
            .I(N__27003));
    InMux I__4462 (
            .O(N__27003),
            .I(N__27000));
    LocalMux I__4461 (
            .O(N__27000),
            .I(N__26997));
    Odrv12 I__4460 (
            .O(N__26997),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ));
    InMux I__4459 (
            .O(N__26994),
            .I(N__26991));
    LocalMux I__4458 (
            .O(N__26991),
            .I(\current_shift_inst.control_input_1_axb_23 ));
    InMux I__4457 (
            .O(N__26988),
            .I(\current_shift_inst.un38_control_input_0_cry_28 ));
    InMux I__4456 (
            .O(N__26985),
            .I(N__26982));
    LocalMux I__4455 (
            .O(N__26982),
            .I(N__26979));
    Span4Mux_h I__4454 (
            .O(N__26979),
            .I(N__26976));
    Odrv4 I__4453 (
            .O(N__26976),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ));
    CascadeMux I__4452 (
            .O(N__26973),
            .I(N__26970));
    InMux I__4451 (
            .O(N__26970),
            .I(N__26966));
    InMux I__4450 (
            .O(N__26969),
            .I(N__26963));
    LocalMux I__4449 (
            .O(N__26966),
            .I(N__26960));
    LocalMux I__4448 (
            .O(N__26963),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ));
    Odrv12 I__4447 (
            .O(N__26960),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ));
    InMux I__4446 (
            .O(N__26955),
            .I(N__26952));
    LocalMux I__4445 (
            .O(N__26952),
            .I(\current_shift_inst.control_input_1_axb_24 ));
    InMux I__4444 (
            .O(N__26949),
            .I(\current_shift_inst.un38_control_input_0_cry_29 ));
    InMux I__4443 (
            .O(N__26946),
            .I(N__26943));
    LocalMux I__4442 (
            .O(N__26943),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    InMux I__4441 (
            .O(N__26940),
            .I(bfn_9_15_0_));
    InMux I__4440 (
            .O(N__26937),
            .I(N__26934));
    LocalMux I__4439 (
            .O(N__26934),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    InMux I__4438 (
            .O(N__26931),
            .I(\current_shift_inst.un38_control_input_0_cry_15 ));
    InMux I__4437 (
            .O(N__26928),
            .I(N__26925));
    LocalMux I__4436 (
            .O(N__26925),
            .I(\current_shift_inst.control_input_1_axb_11 ));
    InMux I__4435 (
            .O(N__26922),
            .I(\current_shift_inst.un38_control_input_0_cry_16 ));
    InMux I__4434 (
            .O(N__26919),
            .I(N__26916));
    LocalMux I__4433 (
            .O(N__26916),
            .I(N__26913));
    Span4Mux_v I__4432 (
            .O(N__26913),
            .I(N__26910));
    Odrv4 I__4431 (
            .O(N__26910),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ));
    InMux I__4430 (
            .O(N__26907),
            .I(N__26904));
    LocalMux I__4429 (
            .O(N__26904),
            .I(\current_shift_inst.control_input_1_axb_12 ));
    InMux I__4428 (
            .O(N__26901),
            .I(\current_shift_inst.un38_control_input_0_cry_17 ));
    InMux I__4427 (
            .O(N__26898),
            .I(N__26895));
    LocalMux I__4426 (
            .O(N__26895),
            .I(N__26892));
    Odrv4 I__4425 (
            .O(N__26892),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ));
    CascadeMux I__4424 (
            .O(N__26889),
            .I(N__26886));
    InMux I__4423 (
            .O(N__26886),
            .I(N__26883));
    LocalMux I__4422 (
            .O(N__26883),
            .I(N__26880));
    Span4Mux_v I__4421 (
            .O(N__26880),
            .I(N__26877));
    Odrv4 I__4420 (
            .O(N__26877),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ));
    InMux I__4419 (
            .O(N__26874),
            .I(N__26871));
    LocalMux I__4418 (
            .O(N__26871),
            .I(\current_shift_inst.control_input_1_axb_13 ));
    InMux I__4417 (
            .O(N__26868),
            .I(\current_shift_inst.un38_control_input_0_cry_18 ));
    InMux I__4416 (
            .O(N__26865),
            .I(N__26862));
    LocalMux I__4415 (
            .O(N__26862),
            .I(N__26859));
    Odrv4 I__4414 (
            .O(N__26859),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ));
    CascadeMux I__4413 (
            .O(N__26856),
            .I(N__26853));
    InMux I__4412 (
            .O(N__26853),
            .I(N__26850));
    LocalMux I__4411 (
            .O(N__26850),
            .I(N__26847));
    Odrv12 I__4410 (
            .O(N__26847),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ));
    InMux I__4409 (
            .O(N__26844),
            .I(N__26841));
    LocalMux I__4408 (
            .O(N__26841),
            .I(\current_shift_inst.control_input_1_axb_14 ));
    InMux I__4407 (
            .O(N__26838),
            .I(\current_shift_inst.un38_control_input_0_cry_19 ));
    InMux I__4406 (
            .O(N__26835),
            .I(N__26832));
    LocalMux I__4405 (
            .O(N__26832),
            .I(N__26829));
    Odrv4 I__4404 (
            .O(N__26829),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ));
    CascadeMux I__4403 (
            .O(N__26826),
            .I(N__26823));
    InMux I__4402 (
            .O(N__26823),
            .I(N__26820));
    LocalMux I__4401 (
            .O(N__26820),
            .I(N__26817));
    Odrv12 I__4400 (
            .O(N__26817),
            .I(\current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ));
    InMux I__4399 (
            .O(N__26814),
            .I(N__26811));
    LocalMux I__4398 (
            .O(N__26811),
            .I(\current_shift_inst.control_input_1_axb_15 ));
    InMux I__4397 (
            .O(N__26808),
            .I(\current_shift_inst.un38_control_input_0_cry_20 ));
    InMux I__4396 (
            .O(N__26805),
            .I(N__26802));
    LocalMux I__4395 (
            .O(N__26802),
            .I(N__26799));
    Odrv4 I__4394 (
            .O(N__26799),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ));
    CascadeMux I__4393 (
            .O(N__26796),
            .I(N__26793));
    InMux I__4392 (
            .O(N__26793),
            .I(N__26790));
    LocalMux I__4391 (
            .O(N__26790),
            .I(N__26787));
    Odrv4 I__4390 (
            .O(N__26787),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ));
    InMux I__4389 (
            .O(N__26784),
            .I(N__26781));
    LocalMux I__4388 (
            .O(N__26781),
            .I(\current_shift_inst.control_input_1_axb_16 ));
    InMux I__4387 (
            .O(N__26778),
            .I(\current_shift_inst.un38_control_input_0_cry_21 ));
    InMux I__4386 (
            .O(N__26775),
            .I(bfn_9_14_0_));
    InMux I__4385 (
            .O(N__26772),
            .I(N__26769));
    LocalMux I__4384 (
            .O(N__26769),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__4383 (
            .O(N__26766),
            .I(\current_shift_inst.un38_control_input_0_cry_7 ));
    InMux I__4382 (
            .O(N__26763),
            .I(N__26760));
    LocalMux I__4381 (
            .O(N__26760),
            .I(N__26757));
    Odrv4 I__4380 (
            .O(N__26757),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ));
    InMux I__4379 (
            .O(N__26754),
            .I(N__26751));
    LocalMux I__4378 (
            .O(N__26751),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    InMux I__4377 (
            .O(N__26748),
            .I(\current_shift_inst.un38_control_input_0_cry_8 ));
    InMux I__4376 (
            .O(N__26745),
            .I(N__26742));
    LocalMux I__4375 (
            .O(N__26742),
            .I(N__26739));
    Odrv4 I__4374 (
            .O(N__26739),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ));
    CascadeMux I__4373 (
            .O(N__26736),
            .I(N__26733));
    InMux I__4372 (
            .O(N__26733),
            .I(N__26730));
    LocalMux I__4371 (
            .O(N__26730),
            .I(N__26727));
    Span4Mux_h I__4370 (
            .O(N__26727),
            .I(N__26724));
    Odrv4 I__4369 (
            .O(N__26724),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ));
    InMux I__4368 (
            .O(N__26721),
            .I(N__26718));
    LocalMux I__4367 (
            .O(N__26718),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__4366 (
            .O(N__26715),
            .I(\current_shift_inst.un38_control_input_0_cry_9 ));
    InMux I__4365 (
            .O(N__26712),
            .I(N__26709));
    LocalMux I__4364 (
            .O(N__26709),
            .I(N__26706));
    Odrv4 I__4363 (
            .O(N__26706),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ));
    CascadeMux I__4362 (
            .O(N__26703),
            .I(N__26700));
    InMux I__4361 (
            .O(N__26700),
            .I(N__26697));
    LocalMux I__4360 (
            .O(N__26697),
            .I(N__26694));
    Span4Mux_h I__4359 (
            .O(N__26694),
            .I(N__26691));
    Odrv4 I__4358 (
            .O(N__26691),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ));
    InMux I__4357 (
            .O(N__26688),
            .I(N__26685));
    LocalMux I__4356 (
            .O(N__26685),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    InMux I__4355 (
            .O(N__26682),
            .I(\current_shift_inst.un38_control_input_0_cry_10 ));
    CascadeMux I__4354 (
            .O(N__26679),
            .I(N__26676));
    InMux I__4353 (
            .O(N__26676),
            .I(N__26673));
    LocalMux I__4352 (
            .O(N__26673),
            .I(N__26670));
    Odrv4 I__4351 (
            .O(N__26670),
            .I(\current_shift_inst.elapsed_time_ns_1_RNILORI_11 ));
    InMux I__4350 (
            .O(N__26667),
            .I(N__26664));
    LocalMux I__4349 (
            .O(N__26664),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    InMux I__4348 (
            .O(N__26661),
            .I(\current_shift_inst.un38_control_input_0_cry_11 ));
    InMux I__4347 (
            .O(N__26658),
            .I(N__26655));
    LocalMux I__4346 (
            .O(N__26655),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__4345 (
            .O(N__26652),
            .I(\current_shift_inst.un38_control_input_0_cry_12 ));
    CascadeMux I__4344 (
            .O(N__26649),
            .I(N__26646));
    InMux I__4343 (
            .O(N__26646),
            .I(N__26643));
    LocalMux I__4342 (
            .O(N__26643),
            .I(N__26640));
    Odrv4 I__4341 (
            .O(N__26640),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ));
    InMux I__4340 (
            .O(N__26637),
            .I(N__26634));
    LocalMux I__4339 (
            .O(N__26634),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    InMux I__4338 (
            .O(N__26631),
            .I(\current_shift_inst.un38_control_input_0_cry_13 ));
    InMux I__4337 (
            .O(N__26628),
            .I(N__26625));
    LocalMux I__4336 (
            .O(N__26625),
            .I(\current_shift_inst.z_i_0_31 ));
    CascadeMux I__4335 (
            .O(N__26622),
            .I(N__26619));
    InMux I__4334 (
            .O(N__26619),
            .I(N__26616));
    LocalMux I__4333 (
            .O(N__26616),
            .I(\current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ));
    InMux I__4332 (
            .O(N__26613),
            .I(N__26610));
    LocalMux I__4331 (
            .O(N__26610),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    InMux I__4330 (
            .O(N__26607),
            .I(\current_shift_inst.un38_control_input_0_cry_5 ));
    InMux I__4329 (
            .O(N__26604),
            .I(N__26601));
    LocalMux I__4328 (
            .O(N__26601),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__4327 (
            .O(N__26598),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ));
    InMux I__4326 (
            .O(N__26595),
            .I(N__26571));
    InMux I__4325 (
            .O(N__26594),
            .I(N__26571));
    InMux I__4324 (
            .O(N__26593),
            .I(N__26571));
    InMux I__4323 (
            .O(N__26592),
            .I(N__26571));
    InMux I__4322 (
            .O(N__26591),
            .I(N__26562));
    InMux I__4321 (
            .O(N__26590),
            .I(N__26562));
    InMux I__4320 (
            .O(N__26589),
            .I(N__26562));
    InMux I__4319 (
            .O(N__26588),
            .I(N__26562));
    InMux I__4318 (
            .O(N__26587),
            .I(N__26553));
    InMux I__4317 (
            .O(N__26586),
            .I(N__26553));
    InMux I__4316 (
            .O(N__26585),
            .I(N__26553));
    InMux I__4315 (
            .O(N__26584),
            .I(N__26553));
    InMux I__4314 (
            .O(N__26583),
            .I(N__26544));
    InMux I__4313 (
            .O(N__26582),
            .I(N__26544));
    InMux I__4312 (
            .O(N__26581),
            .I(N__26544));
    InMux I__4311 (
            .O(N__26580),
            .I(N__26544));
    LocalMux I__4310 (
            .O(N__26571),
            .I(N__26525));
    LocalMux I__4309 (
            .O(N__26562),
            .I(N__26525));
    LocalMux I__4308 (
            .O(N__26553),
            .I(N__26520));
    LocalMux I__4307 (
            .O(N__26544),
            .I(N__26520));
    InMux I__4306 (
            .O(N__26543),
            .I(N__26511));
    InMux I__4305 (
            .O(N__26542),
            .I(N__26511));
    InMux I__4304 (
            .O(N__26541),
            .I(N__26511));
    InMux I__4303 (
            .O(N__26540),
            .I(N__26511));
    InMux I__4302 (
            .O(N__26539),
            .I(N__26502));
    InMux I__4301 (
            .O(N__26538),
            .I(N__26502));
    InMux I__4300 (
            .O(N__26537),
            .I(N__26502));
    InMux I__4299 (
            .O(N__26536),
            .I(N__26502));
    InMux I__4298 (
            .O(N__26535),
            .I(N__26497));
    InMux I__4297 (
            .O(N__26534),
            .I(N__26497));
    InMux I__4296 (
            .O(N__26533),
            .I(N__26488));
    InMux I__4295 (
            .O(N__26532),
            .I(N__26488));
    InMux I__4294 (
            .O(N__26531),
            .I(N__26488));
    InMux I__4293 (
            .O(N__26530),
            .I(N__26488));
    Span4Mux_h I__4292 (
            .O(N__26525),
            .I(N__26485));
    Span4Mux_v I__4291 (
            .O(N__26520),
            .I(N__26482));
    LocalMux I__4290 (
            .O(N__26511),
            .I(\current_shift_inst.timer_phase.running_i ));
    LocalMux I__4289 (
            .O(N__26502),
            .I(\current_shift_inst.timer_phase.running_i ));
    LocalMux I__4288 (
            .O(N__26497),
            .I(\current_shift_inst.timer_phase.running_i ));
    LocalMux I__4287 (
            .O(N__26488),
            .I(\current_shift_inst.timer_phase.running_i ));
    Odrv4 I__4286 (
            .O(N__26485),
            .I(\current_shift_inst.timer_phase.running_i ));
    Odrv4 I__4285 (
            .O(N__26482),
            .I(\current_shift_inst.timer_phase.running_i ));
    InMux I__4284 (
            .O(N__26469),
            .I(N__26466));
    LocalMux I__4283 (
            .O(N__26466),
            .I(N__26463));
    Odrv12 I__4282 (
            .O(N__26463),
            .I(il_min_comp1_c));
    InMux I__4281 (
            .O(N__26460),
            .I(N__26457));
    LocalMux I__4280 (
            .O(N__26457),
            .I(\current_shift_inst.S1_syncZ0Z0 ));
    InMux I__4279 (
            .O(N__26454),
            .I(N__26448));
    InMux I__4278 (
            .O(N__26453),
            .I(N__26448));
    LocalMux I__4277 (
            .O(N__26448),
            .I(\current_shift_inst.S1_syncZ0Z1 ));
    InMux I__4276 (
            .O(N__26445),
            .I(N__26442));
    LocalMux I__4275 (
            .O(N__26442),
            .I(\current_shift_inst.S1_sync_prevZ0 ));
    CascadeMux I__4274 (
            .O(N__26439),
            .I(N__26436));
    InMux I__4273 (
            .O(N__26436),
            .I(N__26432));
    InMux I__4272 (
            .O(N__26435),
            .I(N__26429));
    LocalMux I__4271 (
            .O(N__26432),
            .I(N__26423));
    LocalMux I__4270 (
            .O(N__26429),
            .I(N__26423));
    InMux I__4269 (
            .O(N__26428),
            .I(N__26420));
    Span4Mux_h I__4268 (
            .O(N__26423),
            .I(N__26417));
    LocalMux I__4267 (
            .O(N__26420),
            .I(\current_shift_inst.timer_phase.counterZ0Z_20 ));
    Odrv4 I__4266 (
            .O(N__26417),
            .I(\current_shift_inst.timer_phase.counterZ0Z_20 ));
    InMux I__4265 (
            .O(N__26412),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__4264 (
            .O(N__26409),
            .I(N__26406));
    InMux I__4263 (
            .O(N__26406),
            .I(N__26402));
    InMux I__4262 (
            .O(N__26405),
            .I(N__26399));
    LocalMux I__4261 (
            .O(N__26402),
            .I(N__26393));
    LocalMux I__4260 (
            .O(N__26399),
            .I(N__26393));
    InMux I__4259 (
            .O(N__26398),
            .I(N__26390));
    Span4Mux_h I__4258 (
            .O(N__26393),
            .I(N__26387));
    LocalMux I__4257 (
            .O(N__26390),
            .I(\current_shift_inst.timer_phase.counterZ0Z_21 ));
    Odrv4 I__4256 (
            .O(N__26387),
            .I(\current_shift_inst.timer_phase.counterZ0Z_21 ));
    InMux I__4255 (
            .O(N__26382),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ));
    InMux I__4254 (
            .O(N__26379),
            .I(N__26372));
    InMux I__4253 (
            .O(N__26378),
            .I(N__26372));
    InMux I__4252 (
            .O(N__26377),
            .I(N__26369));
    LocalMux I__4251 (
            .O(N__26372),
            .I(N__26366));
    LocalMux I__4250 (
            .O(N__26369),
            .I(\current_shift_inst.timer_phase.counterZ0Z_22 ));
    Odrv4 I__4249 (
            .O(N__26366),
            .I(\current_shift_inst.timer_phase.counterZ0Z_22 ));
    InMux I__4248 (
            .O(N__26361),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ));
    InMux I__4247 (
            .O(N__26358),
            .I(N__26351));
    InMux I__4246 (
            .O(N__26357),
            .I(N__26351));
    InMux I__4245 (
            .O(N__26356),
            .I(N__26348));
    LocalMux I__4244 (
            .O(N__26351),
            .I(N__26345));
    LocalMux I__4243 (
            .O(N__26348),
            .I(\current_shift_inst.timer_phase.counterZ0Z_23 ));
    Odrv4 I__4242 (
            .O(N__26345),
            .I(\current_shift_inst.timer_phase.counterZ0Z_23 ));
    InMux I__4241 (
            .O(N__26340),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__4240 (
            .O(N__26337),
            .I(N__26333));
    InMux I__4239 (
            .O(N__26336),
            .I(N__26329));
    InMux I__4238 (
            .O(N__26333),
            .I(N__26326));
    InMux I__4237 (
            .O(N__26332),
            .I(N__26323));
    LocalMux I__4236 (
            .O(N__26329),
            .I(N__26318));
    LocalMux I__4235 (
            .O(N__26326),
            .I(N__26318));
    LocalMux I__4234 (
            .O(N__26323),
            .I(\current_shift_inst.timer_phase.counterZ0Z_24 ));
    Odrv4 I__4233 (
            .O(N__26318),
            .I(\current_shift_inst.timer_phase.counterZ0Z_24 ));
    InMux I__4232 (
            .O(N__26313),
            .I(bfn_8_20_0_));
    CascadeMux I__4231 (
            .O(N__26310),
            .I(N__26306));
    InMux I__4230 (
            .O(N__26309),
            .I(N__26302));
    InMux I__4229 (
            .O(N__26306),
            .I(N__26299));
    InMux I__4228 (
            .O(N__26305),
            .I(N__26296));
    LocalMux I__4227 (
            .O(N__26302),
            .I(N__26291));
    LocalMux I__4226 (
            .O(N__26299),
            .I(N__26291));
    LocalMux I__4225 (
            .O(N__26296),
            .I(\current_shift_inst.timer_phase.counterZ0Z_25 ));
    Odrv4 I__4224 (
            .O(N__26291),
            .I(\current_shift_inst.timer_phase.counterZ0Z_25 ));
    InMux I__4223 (
            .O(N__26286),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ));
    InMux I__4222 (
            .O(N__26283),
            .I(N__26280));
    LocalMux I__4221 (
            .O(N__26280),
            .I(N__26276));
    InMux I__4220 (
            .O(N__26279),
            .I(N__26273));
    Span4Mux_h I__4219 (
            .O(N__26276),
            .I(N__26270));
    LocalMux I__4218 (
            .O(N__26273),
            .I(\current_shift_inst.timer_phase.counterZ0Z_28 ));
    Odrv4 I__4217 (
            .O(N__26270),
            .I(\current_shift_inst.timer_phase.counterZ0Z_28 ));
    CascadeMux I__4216 (
            .O(N__26265),
            .I(N__26261));
    CascadeMux I__4215 (
            .O(N__26264),
            .I(N__26258));
    InMux I__4214 (
            .O(N__26261),
            .I(N__26252));
    InMux I__4213 (
            .O(N__26258),
            .I(N__26252));
    InMux I__4212 (
            .O(N__26257),
            .I(N__26249));
    LocalMux I__4211 (
            .O(N__26252),
            .I(N__26246));
    LocalMux I__4210 (
            .O(N__26249),
            .I(\current_shift_inst.timer_phase.counterZ0Z_26 ));
    Odrv4 I__4209 (
            .O(N__26246),
            .I(\current_shift_inst.timer_phase.counterZ0Z_26 ));
    InMux I__4208 (
            .O(N__26241),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ));
    InMux I__4207 (
            .O(N__26238),
            .I(N__26235));
    LocalMux I__4206 (
            .O(N__26235),
            .I(N__26231));
    InMux I__4205 (
            .O(N__26234),
            .I(N__26228));
    Span4Mux_h I__4204 (
            .O(N__26231),
            .I(N__26225));
    LocalMux I__4203 (
            .O(N__26228),
            .I(\current_shift_inst.timer_phase.counterZ0Z_29 ));
    Odrv4 I__4202 (
            .O(N__26225),
            .I(\current_shift_inst.timer_phase.counterZ0Z_29 ));
    CascadeMux I__4201 (
            .O(N__26220),
            .I(N__26216));
    CascadeMux I__4200 (
            .O(N__26219),
            .I(N__26213));
    InMux I__4199 (
            .O(N__26216),
            .I(N__26207));
    InMux I__4198 (
            .O(N__26213),
            .I(N__26207));
    InMux I__4197 (
            .O(N__26212),
            .I(N__26204));
    LocalMux I__4196 (
            .O(N__26207),
            .I(N__26201));
    LocalMux I__4195 (
            .O(N__26204),
            .I(\current_shift_inst.timer_phase.counterZ0Z_27 ));
    Odrv4 I__4194 (
            .O(N__26201),
            .I(\current_shift_inst.timer_phase.counterZ0Z_27 ));
    InMux I__4193 (
            .O(N__26196),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ));
    CascadeMux I__4192 (
            .O(N__26193),
            .I(N__26190));
    InMux I__4191 (
            .O(N__26190),
            .I(N__26186));
    InMux I__4190 (
            .O(N__26189),
            .I(N__26183));
    LocalMux I__4189 (
            .O(N__26186),
            .I(N__26177));
    LocalMux I__4188 (
            .O(N__26183),
            .I(N__26177));
    InMux I__4187 (
            .O(N__26182),
            .I(N__26174));
    Span4Mux_h I__4186 (
            .O(N__26177),
            .I(N__26171));
    LocalMux I__4185 (
            .O(N__26174),
            .I(\current_shift_inst.timer_phase.counterZ0Z_12 ));
    Odrv4 I__4184 (
            .O(N__26171),
            .I(\current_shift_inst.timer_phase.counterZ0Z_12 ));
    InMux I__4183 (
            .O(N__26166),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__4182 (
            .O(N__26163),
            .I(N__26160));
    InMux I__4181 (
            .O(N__26160),
            .I(N__26156));
    InMux I__4180 (
            .O(N__26159),
            .I(N__26153));
    LocalMux I__4179 (
            .O(N__26156),
            .I(N__26147));
    LocalMux I__4178 (
            .O(N__26153),
            .I(N__26147));
    InMux I__4177 (
            .O(N__26152),
            .I(N__26144));
    Span4Mux_h I__4176 (
            .O(N__26147),
            .I(N__26141));
    LocalMux I__4175 (
            .O(N__26144),
            .I(\current_shift_inst.timer_phase.counterZ0Z_13 ));
    Odrv4 I__4174 (
            .O(N__26141),
            .I(\current_shift_inst.timer_phase.counterZ0Z_13 ));
    InMux I__4173 (
            .O(N__26136),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ));
    InMux I__4172 (
            .O(N__26133),
            .I(N__26126));
    InMux I__4171 (
            .O(N__26132),
            .I(N__26126));
    InMux I__4170 (
            .O(N__26131),
            .I(N__26123));
    LocalMux I__4169 (
            .O(N__26126),
            .I(N__26120));
    LocalMux I__4168 (
            .O(N__26123),
            .I(\current_shift_inst.timer_phase.counterZ0Z_14 ));
    Odrv4 I__4167 (
            .O(N__26120),
            .I(\current_shift_inst.timer_phase.counterZ0Z_14 ));
    InMux I__4166 (
            .O(N__26115),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ));
    InMux I__4165 (
            .O(N__26112),
            .I(N__26105));
    InMux I__4164 (
            .O(N__26111),
            .I(N__26105));
    InMux I__4163 (
            .O(N__26110),
            .I(N__26102));
    LocalMux I__4162 (
            .O(N__26105),
            .I(N__26099));
    LocalMux I__4161 (
            .O(N__26102),
            .I(\current_shift_inst.timer_phase.counterZ0Z_15 ));
    Odrv4 I__4160 (
            .O(N__26099),
            .I(\current_shift_inst.timer_phase.counterZ0Z_15 ));
    InMux I__4159 (
            .O(N__26094),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__4158 (
            .O(N__26091),
            .I(N__26087));
    InMux I__4157 (
            .O(N__26090),
            .I(N__26083));
    InMux I__4156 (
            .O(N__26087),
            .I(N__26080));
    InMux I__4155 (
            .O(N__26086),
            .I(N__26077));
    LocalMux I__4154 (
            .O(N__26083),
            .I(N__26072));
    LocalMux I__4153 (
            .O(N__26080),
            .I(N__26072));
    LocalMux I__4152 (
            .O(N__26077),
            .I(\current_shift_inst.timer_phase.counterZ0Z_16 ));
    Odrv4 I__4151 (
            .O(N__26072),
            .I(\current_shift_inst.timer_phase.counterZ0Z_16 ));
    InMux I__4150 (
            .O(N__26067),
            .I(bfn_8_19_0_));
    CascadeMux I__4149 (
            .O(N__26064),
            .I(N__26060));
    InMux I__4148 (
            .O(N__26063),
            .I(N__26056));
    InMux I__4147 (
            .O(N__26060),
            .I(N__26053));
    InMux I__4146 (
            .O(N__26059),
            .I(N__26050));
    LocalMux I__4145 (
            .O(N__26056),
            .I(N__26045));
    LocalMux I__4144 (
            .O(N__26053),
            .I(N__26045));
    LocalMux I__4143 (
            .O(N__26050),
            .I(\current_shift_inst.timer_phase.counterZ0Z_17 ));
    Odrv4 I__4142 (
            .O(N__26045),
            .I(\current_shift_inst.timer_phase.counterZ0Z_17 ));
    InMux I__4141 (
            .O(N__26040),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__4140 (
            .O(N__26037),
            .I(N__26033));
    CascadeMux I__4139 (
            .O(N__26036),
            .I(N__26030));
    InMux I__4138 (
            .O(N__26033),
            .I(N__26024));
    InMux I__4137 (
            .O(N__26030),
            .I(N__26024));
    InMux I__4136 (
            .O(N__26029),
            .I(N__26021));
    LocalMux I__4135 (
            .O(N__26024),
            .I(N__26018));
    LocalMux I__4134 (
            .O(N__26021),
            .I(\current_shift_inst.timer_phase.counterZ0Z_18 ));
    Odrv4 I__4133 (
            .O(N__26018),
            .I(\current_shift_inst.timer_phase.counterZ0Z_18 ));
    InMux I__4132 (
            .O(N__26013),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__4131 (
            .O(N__26010),
            .I(N__26006));
    CascadeMux I__4130 (
            .O(N__26009),
            .I(N__26003));
    InMux I__4129 (
            .O(N__26006),
            .I(N__25997));
    InMux I__4128 (
            .O(N__26003),
            .I(N__25997));
    InMux I__4127 (
            .O(N__26002),
            .I(N__25994));
    LocalMux I__4126 (
            .O(N__25997),
            .I(N__25991));
    LocalMux I__4125 (
            .O(N__25994),
            .I(\current_shift_inst.timer_phase.counterZ0Z_19 ));
    Odrv4 I__4124 (
            .O(N__25991),
            .I(\current_shift_inst.timer_phase.counterZ0Z_19 ));
    InMux I__4123 (
            .O(N__25986),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__4122 (
            .O(N__25983),
            .I(N__25979));
    CascadeMux I__4121 (
            .O(N__25982),
            .I(N__25976));
    InMux I__4120 (
            .O(N__25979),
            .I(N__25970));
    InMux I__4119 (
            .O(N__25976),
            .I(N__25970));
    InMux I__4118 (
            .O(N__25975),
            .I(N__25967));
    LocalMux I__4117 (
            .O(N__25970),
            .I(N__25964));
    LocalMux I__4116 (
            .O(N__25967),
            .I(\current_shift_inst.timer_phase.counterZ0Z_3 ));
    Odrv4 I__4115 (
            .O(N__25964),
            .I(\current_shift_inst.timer_phase.counterZ0Z_3 ));
    InMux I__4114 (
            .O(N__25959),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ));
    InMux I__4113 (
            .O(N__25956),
            .I(N__25950));
    InMux I__4112 (
            .O(N__25955),
            .I(N__25950));
    LocalMux I__4111 (
            .O(N__25950),
            .I(N__25946));
    InMux I__4110 (
            .O(N__25949),
            .I(N__25943));
    Span4Mux_h I__4109 (
            .O(N__25946),
            .I(N__25940));
    LocalMux I__4108 (
            .O(N__25943),
            .I(\current_shift_inst.timer_phase.counterZ0Z_4 ));
    Odrv4 I__4107 (
            .O(N__25940),
            .I(\current_shift_inst.timer_phase.counterZ0Z_4 ));
    InMux I__4106 (
            .O(N__25935),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ));
    InMux I__4105 (
            .O(N__25932),
            .I(N__25925));
    InMux I__4104 (
            .O(N__25931),
            .I(N__25925));
    InMux I__4103 (
            .O(N__25930),
            .I(N__25922));
    LocalMux I__4102 (
            .O(N__25925),
            .I(N__25919));
    LocalMux I__4101 (
            .O(N__25922),
            .I(\current_shift_inst.timer_phase.counterZ0Z_5 ));
    Odrv4 I__4100 (
            .O(N__25919),
            .I(\current_shift_inst.timer_phase.counterZ0Z_5 ));
    InMux I__4099 (
            .O(N__25914),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__4098 (
            .O(N__25911),
            .I(N__25907));
    CascadeMux I__4097 (
            .O(N__25910),
            .I(N__25904));
    InMux I__4096 (
            .O(N__25907),
            .I(N__25899));
    InMux I__4095 (
            .O(N__25904),
            .I(N__25899));
    LocalMux I__4094 (
            .O(N__25899),
            .I(N__25895));
    InMux I__4093 (
            .O(N__25898),
            .I(N__25892));
    Span4Mux_h I__4092 (
            .O(N__25895),
            .I(N__25889));
    LocalMux I__4091 (
            .O(N__25892),
            .I(\current_shift_inst.timer_phase.counterZ0Z_6 ));
    Odrv4 I__4090 (
            .O(N__25889),
            .I(\current_shift_inst.timer_phase.counterZ0Z_6 ));
    InMux I__4089 (
            .O(N__25884),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__4088 (
            .O(N__25881),
            .I(N__25877));
    CascadeMux I__4087 (
            .O(N__25880),
            .I(N__25874));
    InMux I__4086 (
            .O(N__25877),
            .I(N__25869));
    InMux I__4085 (
            .O(N__25874),
            .I(N__25869));
    LocalMux I__4084 (
            .O(N__25869),
            .I(N__25865));
    InMux I__4083 (
            .O(N__25868),
            .I(N__25862));
    Span4Mux_h I__4082 (
            .O(N__25865),
            .I(N__25859));
    LocalMux I__4081 (
            .O(N__25862),
            .I(\current_shift_inst.timer_phase.counterZ0Z_7 ));
    Odrv4 I__4080 (
            .O(N__25859),
            .I(\current_shift_inst.timer_phase.counterZ0Z_7 ));
    InMux I__4079 (
            .O(N__25854),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ));
    InMux I__4078 (
            .O(N__25851),
            .I(N__25847));
    InMux I__4077 (
            .O(N__25850),
            .I(N__25844));
    LocalMux I__4076 (
            .O(N__25847),
            .I(N__25840));
    LocalMux I__4075 (
            .O(N__25844),
            .I(N__25837));
    InMux I__4074 (
            .O(N__25843),
            .I(N__25834));
    Span4Mux_h I__4073 (
            .O(N__25840),
            .I(N__25831));
    Odrv4 I__4072 (
            .O(N__25837),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    LocalMux I__4071 (
            .O(N__25834),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    Odrv4 I__4070 (
            .O(N__25831),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    InMux I__4069 (
            .O(N__25824),
            .I(bfn_8_18_0_));
    InMux I__4068 (
            .O(N__25821),
            .I(N__25817));
    InMux I__4067 (
            .O(N__25820),
            .I(N__25814));
    LocalMux I__4066 (
            .O(N__25817),
            .I(N__25810));
    LocalMux I__4065 (
            .O(N__25814),
            .I(N__25807));
    InMux I__4064 (
            .O(N__25813),
            .I(N__25804));
    Span4Mux_h I__4063 (
            .O(N__25810),
            .I(N__25801));
    Odrv4 I__4062 (
            .O(N__25807),
            .I(\current_shift_inst.timer_phase.counterZ0Z_9 ));
    LocalMux I__4061 (
            .O(N__25804),
            .I(\current_shift_inst.timer_phase.counterZ0Z_9 ));
    Odrv4 I__4060 (
            .O(N__25801),
            .I(\current_shift_inst.timer_phase.counterZ0Z_9 ));
    InMux I__4059 (
            .O(N__25794),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__4058 (
            .O(N__25791),
            .I(N__25787));
    CascadeMux I__4057 (
            .O(N__25790),
            .I(N__25784));
    InMux I__4056 (
            .O(N__25787),
            .I(N__25778));
    InMux I__4055 (
            .O(N__25784),
            .I(N__25778));
    InMux I__4054 (
            .O(N__25783),
            .I(N__25775));
    LocalMux I__4053 (
            .O(N__25778),
            .I(N__25772));
    LocalMux I__4052 (
            .O(N__25775),
            .I(\current_shift_inst.timer_phase.counterZ0Z_10 ));
    Odrv4 I__4051 (
            .O(N__25772),
            .I(\current_shift_inst.timer_phase.counterZ0Z_10 ));
    InMux I__4050 (
            .O(N__25767),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__4049 (
            .O(N__25764),
            .I(N__25760));
    CascadeMux I__4048 (
            .O(N__25763),
            .I(N__25757));
    InMux I__4047 (
            .O(N__25760),
            .I(N__25751));
    InMux I__4046 (
            .O(N__25757),
            .I(N__25751));
    InMux I__4045 (
            .O(N__25756),
            .I(N__25748));
    LocalMux I__4044 (
            .O(N__25751),
            .I(N__25745));
    LocalMux I__4043 (
            .O(N__25748),
            .I(\current_shift_inst.timer_phase.counterZ0Z_11 ));
    Odrv4 I__4042 (
            .O(N__25745),
            .I(\current_shift_inst.timer_phase.counterZ0Z_11 ));
    InMux I__4041 (
            .O(N__25740),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__4040 (
            .O(N__25737),
            .I(N__25734));
    InMux I__4039 (
            .O(N__25734),
            .I(N__25730));
    InMux I__4038 (
            .O(N__25733),
            .I(N__25727));
    LocalMux I__4037 (
            .O(N__25730),
            .I(N__25724));
    LocalMux I__4036 (
            .O(N__25727),
            .I(N__25721));
    Span4Mux_v I__4035 (
            .O(N__25724),
            .I(N__25718));
    Odrv4 I__4034 (
            .O(N__25721),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    Odrv4 I__4033 (
            .O(N__25718),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    InMux I__4032 (
            .O(N__25713),
            .I(\current_shift_inst.control_input_1_cry_20 ));
    CascadeMux I__4031 (
            .O(N__25710),
            .I(N__25706));
    InMux I__4030 (
            .O(N__25709),
            .I(N__25703));
    InMux I__4029 (
            .O(N__25706),
            .I(N__25700));
    LocalMux I__4028 (
            .O(N__25703),
            .I(N__25697));
    LocalMux I__4027 (
            .O(N__25700),
            .I(N__25694));
    Span4Mux_h I__4026 (
            .O(N__25697),
            .I(N__25689));
    Span4Mux_h I__4025 (
            .O(N__25694),
            .I(N__25689));
    Odrv4 I__4024 (
            .O(N__25689),
            .I(\current_shift_inst.control_inputZ0Z_22 ));
    InMux I__4023 (
            .O(N__25686),
            .I(\current_shift_inst.control_input_1_cry_21 ));
    CascadeMux I__4022 (
            .O(N__25683),
            .I(N__25679));
    InMux I__4021 (
            .O(N__25682),
            .I(N__25676));
    InMux I__4020 (
            .O(N__25679),
            .I(N__25673));
    LocalMux I__4019 (
            .O(N__25676),
            .I(N__25670));
    LocalMux I__4018 (
            .O(N__25673),
            .I(N__25667));
    Span4Mux_h I__4017 (
            .O(N__25670),
            .I(N__25662));
    Span4Mux_h I__4016 (
            .O(N__25667),
            .I(N__25662));
    Odrv4 I__4015 (
            .O(N__25662),
            .I(\current_shift_inst.control_inputZ0Z_23 ));
    InMux I__4014 (
            .O(N__25659),
            .I(\current_shift_inst.control_input_1_cry_22 ));
    CascadeMux I__4013 (
            .O(N__25656),
            .I(N__25653));
    InMux I__4012 (
            .O(N__25653),
            .I(N__25649));
    InMux I__4011 (
            .O(N__25652),
            .I(N__25646));
    LocalMux I__4010 (
            .O(N__25649),
            .I(N__25643));
    LocalMux I__4009 (
            .O(N__25646),
            .I(N__25640));
    Span4Mux_h I__4008 (
            .O(N__25643),
            .I(N__25637));
    Odrv12 I__4007 (
            .O(N__25640),
            .I(\current_shift_inst.control_inputZ0Z_24 ));
    Odrv4 I__4006 (
            .O(N__25637),
            .I(\current_shift_inst.control_inputZ0Z_24 ));
    InMux I__4005 (
            .O(N__25632),
            .I(bfn_8_16_0_));
    InMux I__4004 (
            .O(N__25629),
            .I(\current_shift_inst.control_input_1_cry_24 ));
    InMux I__4003 (
            .O(N__25626),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__4002 (
            .O(N__25623),
            .I(N__25619));
    CascadeMux I__4001 (
            .O(N__25622),
            .I(N__25616));
    InMux I__4000 (
            .O(N__25619),
            .I(N__25610));
    InMux I__3999 (
            .O(N__25616),
            .I(N__25610));
    InMux I__3998 (
            .O(N__25615),
            .I(N__25607));
    LocalMux I__3997 (
            .O(N__25610),
            .I(N__25604));
    LocalMux I__3996 (
            .O(N__25607),
            .I(\current_shift_inst.timer_phase.counterZ0Z_2 ));
    Odrv4 I__3995 (
            .O(N__25604),
            .I(\current_shift_inst.timer_phase.counterZ0Z_2 ));
    InMux I__3994 (
            .O(N__25599),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ));
    InMux I__3993 (
            .O(N__25596),
            .I(N__25592));
    InMux I__3992 (
            .O(N__25595),
            .I(N__25589));
    LocalMux I__3991 (
            .O(N__25592),
            .I(N__25584));
    LocalMux I__3990 (
            .O(N__25589),
            .I(N__25584));
    Span4Mux_v I__3989 (
            .O(N__25584),
            .I(N__25581));
    Odrv4 I__3988 (
            .O(N__25581),
            .I(\current_shift_inst.control_inputZ0Z_12 ));
    InMux I__3987 (
            .O(N__25578),
            .I(\current_shift_inst.control_input_1_cry_11 ));
    CascadeMux I__3986 (
            .O(N__25575),
            .I(N__25571));
    InMux I__3985 (
            .O(N__25574),
            .I(N__25568));
    InMux I__3984 (
            .O(N__25571),
            .I(N__25565));
    LocalMux I__3983 (
            .O(N__25568),
            .I(N__25560));
    LocalMux I__3982 (
            .O(N__25565),
            .I(N__25560));
    Span4Mux_v I__3981 (
            .O(N__25560),
            .I(N__25557));
    Odrv4 I__3980 (
            .O(N__25557),
            .I(\current_shift_inst.control_inputZ0Z_13 ));
    InMux I__3979 (
            .O(N__25554),
            .I(\current_shift_inst.control_input_1_cry_12 ));
    CascadeMux I__3978 (
            .O(N__25551),
            .I(N__25547));
    InMux I__3977 (
            .O(N__25550),
            .I(N__25544));
    InMux I__3976 (
            .O(N__25547),
            .I(N__25541));
    LocalMux I__3975 (
            .O(N__25544),
            .I(N__25536));
    LocalMux I__3974 (
            .O(N__25541),
            .I(N__25536));
    Span4Mux_v I__3973 (
            .O(N__25536),
            .I(N__25533));
    Odrv4 I__3972 (
            .O(N__25533),
            .I(\current_shift_inst.control_inputZ0Z_14 ));
    InMux I__3971 (
            .O(N__25530),
            .I(\current_shift_inst.control_input_1_cry_13 ));
    CascadeMux I__3970 (
            .O(N__25527),
            .I(N__25523));
    InMux I__3969 (
            .O(N__25526),
            .I(N__25520));
    InMux I__3968 (
            .O(N__25523),
            .I(N__25517));
    LocalMux I__3967 (
            .O(N__25520),
            .I(N__25512));
    LocalMux I__3966 (
            .O(N__25517),
            .I(N__25512));
    Span4Mux_v I__3965 (
            .O(N__25512),
            .I(N__25509));
    Odrv4 I__3964 (
            .O(N__25509),
            .I(\current_shift_inst.control_inputZ0Z_15 ));
    InMux I__3963 (
            .O(N__25506),
            .I(\current_shift_inst.control_input_1_cry_14 ));
    CascadeMux I__3962 (
            .O(N__25503),
            .I(N__25500));
    InMux I__3961 (
            .O(N__25500),
            .I(N__25496));
    InMux I__3960 (
            .O(N__25499),
            .I(N__25493));
    LocalMux I__3959 (
            .O(N__25496),
            .I(N__25490));
    LocalMux I__3958 (
            .O(N__25493),
            .I(N__25487));
    Span4Mux_h I__3957 (
            .O(N__25490),
            .I(N__25484));
    Odrv12 I__3956 (
            .O(N__25487),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    Odrv4 I__3955 (
            .O(N__25484),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    InMux I__3954 (
            .O(N__25479),
            .I(bfn_8_15_0_));
    CascadeMux I__3953 (
            .O(N__25476),
            .I(N__25473));
    InMux I__3952 (
            .O(N__25473),
            .I(N__25469));
    InMux I__3951 (
            .O(N__25472),
            .I(N__25466));
    LocalMux I__3950 (
            .O(N__25469),
            .I(N__25463));
    LocalMux I__3949 (
            .O(N__25466),
            .I(N__25460));
    Span12Mux_s8_h I__3948 (
            .O(N__25463),
            .I(N__25457));
    Odrv12 I__3947 (
            .O(N__25460),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    Odrv12 I__3946 (
            .O(N__25457),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    InMux I__3945 (
            .O(N__25452),
            .I(\current_shift_inst.control_input_1_cry_16 ));
    CascadeMux I__3944 (
            .O(N__25449),
            .I(N__25446));
    InMux I__3943 (
            .O(N__25446),
            .I(N__25443));
    LocalMux I__3942 (
            .O(N__25443),
            .I(N__25439));
    InMux I__3941 (
            .O(N__25442),
            .I(N__25436));
    Span4Mux_v I__3940 (
            .O(N__25439),
            .I(N__25433));
    LocalMux I__3939 (
            .O(N__25436),
            .I(N__25430));
    Span4Mux_h I__3938 (
            .O(N__25433),
            .I(N__25427));
    Odrv12 I__3937 (
            .O(N__25430),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    Odrv4 I__3936 (
            .O(N__25427),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    InMux I__3935 (
            .O(N__25422),
            .I(\current_shift_inst.control_input_1_cry_17 ));
    CascadeMux I__3934 (
            .O(N__25419),
            .I(N__25416));
    InMux I__3933 (
            .O(N__25416),
            .I(N__25412));
    InMux I__3932 (
            .O(N__25415),
            .I(N__25409));
    LocalMux I__3931 (
            .O(N__25412),
            .I(N__25406));
    LocalMux I__3930 (
            .O(N__25409),
            .I(N__25403));
    Span4Mux_h I__3929 (
            .O(N__25406),
            .I(N__25400));
    Odrv4 I__3928 (
            .O(N__25403),
            .I(\current_shift_inst.control_inputZ0Z_19 ));
    Odrv4 I__3927 (
            .O(N__25400),
            .I(\current_shift_inst.control_inputZ0Z_19 ));
    InMux I__3926 (
            .O(N__25395),
            .I(\current_shift_inst.control_input_1_cry_18 ));
    CascadeMux I__3925 (
            .O(N__25392),
            .I(N__25389));
    InMux I__3924 (
            .O(N__25389),
            .I(N__25385));
    InMux I__3923 (
            .O(N__25388),
            .I(N__25382));
    LocalMux I__3922 (
            .O(N__25385),
            .I(N__25379));
    LocalMux I__3921 (
            .O(N__25382),
            .I(N__25374));
    Span4Mux_v I__3920 (
            .O(N__25379),
            .I(N__25374));
    Odrv4 I__3919 (
            .O(N__25374),
            .I(\current_shift_inst.control_inputZ0Z_20 ));
    InMux I__3918 (
            .O(N__25371),
            .I(\current_shift_inst.control_input_1_cry_19 ));
    CascadeMux I__3917 (
            .O(N__25368),
            .I(N__25365));
    InMux I__3916 (
            .O(N__25365),
            .I(N__25362));
    LocalMux I__3915 (
            .O(N__25362),
            .I(N__25358));
    InMux I__3914 (
            .O(N__25361),
            .I(N__25355));
    Span4Mux_v I__3913 (
            .O(N__25358),
            .I(N__25352));
    LocalMux I__3912 (
            .O(N__25355),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    Odrv4 I__3911 (
            .O(N__25352),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    InMux I__3910 (
            .O(N__25347),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    InMux I__3909 (
            .O(N__25344),
            .I(N__25340));
    CascadeMux I__3908 (
            .O(N__25343),
            .I(N__25337));
    LocalMux I__3907 (
            .O(N__25340),
            .I(N__25334));
    InMux I__3906 (
            .O(N__25337),
            .I(N__25331));
    Span4Mux_h I__3905 (
            .O(N__25334),
            .I(N__25328));
    LocalMux I__3904 (
            .O(N__25331),
            .I(N__25325));
    Span4Mux_v I__3903 (
            .O(N__25328),
            .I(N__25322));
    Span4Mux_v I__3902 (
            .O(N__25325),
            .I(N__25319));
    Odrv4 I__3901 (
            .O(N__25322),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    Odrv4 I__3900 (
            .O(N__25319),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    InMux I__3899 (
            .O(N__25314),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    CascadeMux I__3898 (
            .O(N__25311),
            .I(N__25307));
    InMux I__3897 (
            .O(N__25310),
            .I(N__25304));
    InMux I__3896 (
            .O(N__25307),
            .I(N__25301));
    LocalMux I__3895 (
            .O(N__25304),
            .I(N__25298));
    LocalMux I__3894 (
            .O(N__25301),
            .I(N__25295));
    Span4Mux_h I__3893 (
            .O(N__25298),
            .I(N__25290));
    Span4Mux_h I__3892 (
            .O(N__25295),
            .I(N__25290));
    Odrv4 I__3891 (
            .O(N__25290),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__3890 (
            .O(N__25287),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    InMux I__3889 (
            .O(N__25284),
            .I(N__25280));
    CascadeMux I__3888 (
            .O(N__25283),
            .I(N__25277));
    LocalMux I__3887 (
            .O(N__25280),
            .I(N__25274));
    InMux I__3886 (
            .O(N__25277),
            .I(N__25271));
    Span4Mux_v I__3885 (
            .O(N__25274),
            .I(N__25266));
    LocalMux I__3884 (
            .O(N__25271),
            .I(N__25266));
    Span4Mux_h I__3883 (
            .O(N__25266),
            .I(N__25263));
    Span4Mux_h I__3882 (
            .O(N__25263),
            .I(N__25260));
    Odrv4 I__3881 (
            .O(N__25260),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    InMux I__3880 (
            .O(N__25257),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    CascadeMux I__3879 (
            .O(N__25254),
            .I(N__25250));
    InMux I__3878 (
            .O(N__25253),
            .I(N__25247));
    InMux I__3877 (
            .O(N__25250),
            .I(N__25244));
    LocalMux I__3876 (
            .O(N__25247),
            .I(N__25241));
    LocalMux I__3875 (
            .O(N__25244),
            .I(N__25238));
    Span4Mux_h I__3874 (
            .O(N__25241),
            .I(N__25235));
    Span4Mux_h I__3873 (
            .O(N__25238),
            .I(N__25232));
    Odrv4 I__3872 (
            .O(N__25235),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    Odrv4 I__3871 (
            .O(N__25232),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__3870 (
            .O(N__25227),
            .I(bfn_8_14_0_));
    InMux I__3869 (
            .O(N__25224),
            .I(N__25220));
    CascadeMux I__3868 (
            .O(N__25223),
            .I(N__25217));
    LocalMux I__3867 (
            .O(N__25220),
            .I(N__25214));
    InMux I__3866 (
            .O(N__25217),
            .I(N__25211));
    Span4Mux_h I__3865 (
            .O(N__25214),
            .I(N__25208));
    LocalMux I__3864 (
            .O(N__25211),
            .I(N__25205));
    Span4Mux_v I__3863 (
            .O(N__25208),
            .I(N__25202));
    Span4Mux_h I__3862 (
            .O(N__25205),
            .I(N__25199));
    Odrv4 I__3861 (
            .O(N__25202),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    Odrv4 I__3860 (
            .O(N__25199),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    InMux I__3859 (
            .O(N__25194),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__3858 (
            .O(N__25191),
            .I(N__25187));
    InMux I__3857 (
            .O(N__25190),
            .I(N__25184));
    LocalMux I__3856 (
            .O(N__25187),
            .I(N__25181));
    LocalMux I__3855 (
            .O(N__25184),
            .I(N__25178));
    Span4Mux_h I__3854 (
            .O(N__25181),
            .I(N__25175));
    Odrv12 I__3853 (
            .O(N__25178),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    Odrv4 I__3852 (
            .O(N__25175),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    InMux I__3851 (
            .O(N__25170),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__3850 (
            .O(N__25167),
            .I(N__25163));
    InMux I__3849 (
            .O(N__25166),
            .I(N__25160));
    LocalMux I__3848 (
            .O(N__25163),
            .I(N__25157));
    LocalMux I__3847 (
            .O(N__25160),
            .I(N__25154));
    Span4Mux_v I__3846 (
            .O(N__25157),
            .I(N__25149));
    Span4Mux_v I__3845 (
            .O(N__25154),
            .I(N__25149));
    Odrv4 I__3844 (
            .O(N__25149),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    InMux I__3843 (
            .O(N__25146),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    InMux I__3842 (
            .O(N__25143),
            .I(N__25140));
    LocalMux I__3841 (
            .O(N__25140),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31 ));
    InMux I__3840 (
            .O(N__25137),
            .I(N__25134));
    LocalMux I__3839 (
            .O(N__25134),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31 ));
    CascadeMux I__3838 (
            .O(N__25131),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31_cascade_ ));
    InMux I__3837 (
            .O(N__25128),
            .I(N__25125));
    LocalMux I__3836 (
            .O(N__25125),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31 ));
    InMux I__3835 (
            .O(N__25122),
            .I(N__25118));
    InMux I__3834 (
            .O(N__25121),
            .I(N__25115));
    LocalMux I__3833 (
            .O(N__25118),
            .I(\current_shift_inst.PI_CTRL.N_47_21 ));
    LocalMux I__3832 (
            .O(N__25115),
            .I(\current_shift_inst.PI_CTRL.N_47_21 ));
    CascadeMux I__3831 (
            .O(N__25110),
            .I(N__25107));
    InMux I__3830 (
            .O(N__25107),
            .I(N__25104));
    LocalMux I__3829 (
            .O(N__25104),
            .I(N__25101));
    Span4Mux_v I__3828 (
            .O(N__25101),
            .I(N__25098));
    Span4Mux_h I__3827 (
            .O(N__25098),
            .I(N__25095));
    Odrv4 I__3826 (
            .O(N__25095),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    CascadeMux I__3825 (
            .O(N__25092),
            .I(N__25089));
    InMux I__3824 (
            .O(N__25089),
            .I(N__25086));
    LocalMux I__3823 (
            .O(N__25086),
            .I(N__25083));
    Span4Mux_h I__3822 (
            .O(N__25083),
            .I(N__25080));
    Odrv4 I__3821 (
            .O(N__25080),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__3820 (
            .O(N__25077),
            .I(N__25073));
    CascadeMux I__3819 (
            .O(N__25076),
            .I(N__25070));
    InMux I__3818 (
            .O(N__25073),
            .I(N__25067));
    InMux I__3817 (
            .O(N__25070),
            .I(N__25064));
    LocalMux I__3816 (
            .O(N__25067),
            .I(N__25061));
    LocalMux I__3815 (
            .O(N__25064),
            .I(N__25058));
    Span4Mux_v I__3814 (
            .O(N__25061),
            .I(N__25053));
    Span4Mux_h I__3813 (
            .O(N__25058),
            .I(N__25050));
    InMux I__3812 (
            .O(N__25057),
            .I(N__25045));
    InMux I__3811 (
            .O(N__25056),
            .I(N__25045));
    Span4Mux_h I__3810 (
            .O(N__25053),
            .I(N__25040));
    Span4Mux_h I__3809 (
            .O(N__25050),
            .I(N__25040));
    LocalMux I__3808 (
            .O(N__25045),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__3807 (
            .O(N__25040),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__3806 (
            .O(N__25035),
            .I(N__25031));
    InMux I__3805 (
            .O(N__25034),
            .I(N__25028));
    LocalMux I__3804 (
            .O(N__25031),
            .I(N__25018));
    LocalMux I__3803 (
            .O(N__25028),
            .I(N__25018));
    InMux I__3802 (
            .O(N__25027),
            .I(N__25009));
    InMux I__3801 (
            .O(N__25026),
            .I(N__25009));
    InMux I__3800 (
            .O(N__25025),
            .I(N__25009));
    InMux I__3799 (
            .O(N__25024),
            .I(N__25009));
    InMux I__3798 (
            .O(N__25023),
            .I(N__25006));
    Span4Mux_v I__3797 (
            .O(N__25018),
            .I(N__24994));
    LocalMux I__3796 (
            .O(N__25009),
            .I(N__24994));
    LocalMux I__3795 (
            .O(N__25006),
            .I(N__24994));
    InMux I__3794 (
            .O(N__25005),
            .I(N__24983));
    InMux I__3793 (
            .O(N__25004),
            .I(N__24983));
    InMux I__3792 (
            .O(N__25003),
            .I(N__24983));
    InMux I__3791 (
            .O(N__25002),
            .I(N__24983));
    InMux I__3790 (
            .O(N__25001),
            .I(N__24983));
    Span4Mux_v I__3789 (
            .O(N__24994),
            .I(N__24964));
    LocalMux I__3788 (
            .O(N__24983),
            .I(N__24964));
    InMux I__3787 (
            .O(N__24982),
            .I(N__24951));
    InMux I__3786 (
            .O(N__24981),
            .I(N__24951));
    InMux I__3785 (
            .O(N__24980),
            .I(N__24951));
    InMux I__3784 (
            .O(N__24979),
            .I(N__24951));
    InMux I__3783 (
            .O(N__24978),
            .I(N__24951));
    InMux I__3782 (
            .O(N__24977),
            .I(N__24951));
    InMux I__3781 (
            .O(N__24976),
            .I(N__24936));
    InMux I__3780 (
            .O(N__24975),
            .I(N__24936));
    InMux I__3779 (
            .O(N__24974),
            .I(N__24936));
    InMux I__3778 (
            .O(N__24973),
            .I(N__24936));
    InMux I__3777 (
            .O(N__24972),
            .I(N__24936));
    InMux I__3776 (
            .O(N__24971),
            .I(N__24936));
    InMux I__3775 (
            .O(N__24970),
            .I(N__24931));
    InMux I__3774 (
            .O(N__24969),
            .I(N__24931));
    Span4Mux_h I__3773 (
            .O(N__24964),
            .I(N__24928));
    LocalMux I__3772 (
            .O(N__24951),
            .I(N__24925));
    InMux I__3771 (
            .O(N__24950),
            .I(N__24920));
    InMux I__3770 (
            .O(N__24949),
            .I(N__24920));
    LocalMux I__3769 (
            .O(N__24936),
            .I(N__24915));
    LocalMux I__3768 (
            .O(N__24931),
            .I(N__24915));
    Odrv4 I__3767 (
            .O(N__24928),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    Odrv12 I__3766 (
            .O(N__24925),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    LocalMux I__3765 (
            .O(N__24920),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    Odrv4 I__3764 (
            .O(N__24915),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    InMux I__3763 (
            .O(N__24906),
            .I(N__24903));
    LocalMux I__3762 (
            .O(N__24903),
            .I(N__24900));
    Odrv4 I__3761 (
            .O(N__24900),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    CascadeMux I__3760 (
            .O(N__24897),
            .I(N__24882));
    CascadeMux I__3759 (
            .O(N__24896),
            .I(N__24879));
    CascadeMux I__3758 (
            .O(N__24895),
            .I(N__24876));
    CascadeMux I__3757 (
            .O(N__24894),
            .I(N__24873));
    CascadeMux I__3756 (
            .O(N__24893),
            .I(N__24868));
    CascadeMux I__3755 (
            .O(N__24892),
            .I(N__24864));
    CascadeMux I__3754 (
            .O(N__24891),
            .I(N__24861));
    CascadeMux I__3753 (
            .O(N__24890),
            .I(N__24858));
    CascadeMux I__3752 (
            .O(N__24889),
            .I(N__24855));
    CascadeMux I__3751 (
            .O(N__24888),
            .I(N__24852));
    CascadeMux I__3750 (
            .O(N__24887),
            .I(N__24847));
    CascadeMux I__3749 (
            .O(N__24886),
            .I(N__24844));
    CascadeMux I__3748 (
            .O(N__24885),
            .I(N__24841));
    InMux I__3747 (
            .O(N__24882),
            .I(N__24829));
    InMux I__3746 (
            .O(N__24879),
            .I(N__24829));
    InMux I__3745 (
            .O(N__24876),
            .I(N__24829));
    InMux I__3744 (
            .O(N__24873),
            .I(N__24829));
    InMux I__3743 (
            .O(N__24872),
            .I(N__24829));
    CascadeMux I__3742 (
            .O(N__24871),
            .I(N__24825));
    InMux I__3741 (
            .O(N__24868),
            .I(N__24815));
    InMux I__3740 (
            .O(N__24867),
            .I(N__24812));
    InMux I__3739 (
            .O(N__24864),
            .I(N__24809));
    InMux I__3738 (
            .O(N__24861),
            .I(N__24804));
    InMux I__3737 (
            .O(N__24858),
            .I(N__24804));
    InMux I__3736 (
            .O(N__24855),
            .I(N__24795));
    InMux I__3735 (
            .O(N__24852),
            .I(N__24795));
    InMux I__3734 (
            .O(N__24851),
            .I(N__24795));
    InMux I__3733 (
            .O(N__24850),
            .I(N__24795));
    InMux I__3732 (
            .O(N__24847),
            .I(N__24786));
    InMux I__3731 (
            .O(N__24844),
            .I(N__24786));
    InMux I__3730 (
            .O(N__24841),
            .I(N__24786));
    InMux I__3729 (
            .O(N__24840),
            .I(N__24786));
    LocalMux I__3728 (
            .O(N__24829),
            .I(N__24783));
    CascadeMux I__3727 (
            .O(N__24828),
            .I(N__24779));
    InMux I__3726 (
            .O(N__24825),
            .I(N__24775));
    InMux I__3725 (
            .O(N__24824),
            .I(N__24770));
    InMux I__3724 (
            .O(N__24823),
            .I(N__24770));
    CascadeMux I__3723 (
            .O(N__24822),
            .I(N__24767));
    CascadeMux I__3722 (
            .O(N__24821),
            .I(N__24763));
    CascadeMux I__3721 (
            .O(N__24820),
            .I(N__24760));
    CascadeMux I__3720 (
            .O(N__24819),
            .I(N__24757));
    CascadeMux I__3719 (
            .O(N__24818),
            .I(N__24754));
    LocalMux I__3718 (
            .O(N__24815),
            .I(N__24749));
    LocalMux I__3717 (
            .O(N__24812),
            .I(N__24746));
    LocalMux I__3716 (
            .O(N__24809),
            .I(N__24739));
    LocalMux I__3715 (
            .O(N__24804),
            .I(N__24739));
    LocalMux I__3714 (
            .O(N__24795),
            .I(N__24739));
    LocalMux I__3713 (
            .O(N__24786),
            .I(N__24734));
    Span4Mux_h I__3712 (
            .O(N__24783),
            .I(N__24734));
    InMux I__3711 (
            .O(N__24782),
            .I(N__24731));
    InMux I__3710 (
            .O(N__24779),
            .I(N__24726));
    InMux I__3709 (
            .O(N__24778),
            .I(N__24726));
    LocalMux I__3708 (
            .O(N__24775),
            .I(N__24723));
    LocalMux I__3707 (
            .O(N__24770),
            .I(N__24720));
    InMux I__3706 (
            .O(N__24767),
            .I(N__24715));
    InMux I__3705 (
            .O(N__24766),
            .I(N__24715));
    InMux I__3704 (
            .O(N__24763),
            .I(N__24702));
    InMux I__3703 (
            .O(N__24760),
            .I(N__24702));
    InMux I__3702 (
            .O(N__24757),
            .I(N__24702));
    InMux I__3701 (
            .O(N__24754),
            .I(N__24702));
    InMux I__3700 (
            .O(N__24753),
            .I(N__24702));
    InMux I__3699 (
            .O(N__24752),
            .I(N__24702));
    Span4Mux_h I__3698 (
            .O(N__24749),
            .I(N__24699));
    Span4Mux_v I__3697 (
            .O(N__24746),
            .I(N__24690));
    Span4Mux_v I__3696 (
            .O(N__24739),
            .I(N__24690));
    Span4Mux_v I__3695 (
            .O(N__24734),
            .I(N__24690));
    LocalMux I__3694 (
            .O(N__24731),
            .I(N__24690));
    LocalMux I__3693 (
            .O(N__24726),
            .I(N__24683));
    Span4Mux_h I__3692 (
            .O(N__24723),
            .I(N__24683));
    Span4Mux_h I__3691 (
            .O(N__24720),
            .I(N__24683));
    LocalMux I__3690 (
            .O(N__24715),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3689 (
            .O(N__24702),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3688 (
            .O(N__24699),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3687 (
            .O(N__24690),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3686 (
            .O(N__24683),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__3685 (
            .O(N__24672),
            .I(N__24667));
    InMux I__3684 (
            .O(N__24671),
            .I(N__24664));
    CascadeMux I__3683 (
            .O(N__24670),
            .I(N__24642));
    LocalMux I__3682 (
            .O(N__24667),
            .I(N__24636));
    LocalMux I__3681 (
            .O(N__24664),
            .I(N__24636));
    InMux I__3680 (
            .O(N__24663),
            .I(N__24627));
    InMux I__3679 (
            .O(N__24662),
            .I(N__24627));
    InMux I__3678 (
            .O(N__24661),
            .I(N__24627));
    InMux I__3677 (
            .O(N__24660),
            .I(N__24627));
    InMux I__3676 (
            .O(N__24659),
            .I(N__24624));
    InMux I__3675 (
            .O(N__24658),
            .I(N__24611));
    InMux I__3674 (
            .O(N__24657),
            .I(N__24611));
    InMux I__3673 (
            .O(N__24656),
            .I(N__24611));
    InMux I__3672 (
            .O(N__24655),
            .I(N__24611));
    InMux I__3671 (
            .O(N__24654),
            .I(N__24611));
    InMux I__3670 (
            .O(N__24653),
            .I(N__24611));
    InMux I__3669 (
            .O(N__24652),
            .I(N__24606));
    InMux I__3668 (
            .O(N__24651),
            .I(N__24606));
    InMux I__3667 (
            .O(N__24650),
            .I(N__24588));
    InMux I__3666 (
            .O(N__24649),
            .I(N__24588));
    InMux I__3665 (
            .O(N__24648),
            .I(N__24588));
    InMux I__3664 (
            .O(N__24647),
            .I(N__24588));
    InMux I__3663 (
            .O(N__24646),
            .I(N__24588));
    InMux I__3662 (
            .O(N__24645),
            .I(N__24588));
    InMux I__3661 (
            .O(N__24642),
            .I(N__24583));
    InMux I__3660 (
            .O(N__24641),
            .I(N__24583));
    Span4Mux_v I__3659 (
            .O(N__24636),
            .I(N__24574));
    LocalMux I__3658 (
            .O(N__24627),
            .I(N__24574));
    LocalMux I__3657 (
            .O(N__24624),
            .I(N__24574));
    LocalMux I__3656 (
            .O(N__24611),
            .I(N__24574));
    LocalMux I__3655 (
            .O(N__24606),
            .I(N__24571));
    InMux I__3654 (
            .O(N__24605),
            .I(N__24560));
    InMux I__3653 (
            .O(N__24604),
            .I(N__24560));
    InMux I__3652 (
            .O(N__24603),
            .I(N__24560));
    InMux I__3651 (
            .O(N__24602),
            .I(N__24560));
    InMux I__3650 (
            .O(N__24601),
            .I(N__24560));
    LocalMux I__3649 (
            .O(N__24588),
            .I(N__24557));
    LocalMux I__3648 (
            .O(N__24583),
            .I(N__24554));
    Span4Mux_v I__3647 (
            .O(N__24574),
            .I(N__24547));
    Span4Mux_v I__3646 (
            .O(N__24571),
            .I(N__24547));
    LocalMux I__3645 (
            .O(N__24560),
            .I(N__24547));
    Odrv12 I__3644 (
            .O(N__24557),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__3643 (
            .O(N__24554),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__3642 (
            .O(N__24547),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    InMux I__3641 (
            .O(N__24540),
            .I(N__24537));
    LocalMux I__3640 (
            .O(N__24537),
            .I(N__24531));
    InMux I__3639 (
            .O(N__24536),
            .I(N__24528));
    InMux I__3638 (
            .O(N__24535),
            .I(N__24523));
    InMux I__3637 (
            .O(N__24534),
            .I(N__24523));
    Span4Mux_v I__3636 (
            .O(N__24531),
            .I(N__24518));
    LocalMux I__3635 (
            .O(N__24528),
            .I(N__24518));
    LocalMux I__3634 (
            .O(N__24523),
            .I(N__24515));
    Odrv4 I__3633 (
            .O(N__24518),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__3632 (
            .O(N__24515),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    CEMux I__3631 (
            .O(N__24510),
            .I(N__24503));
    CEMux I__3630 (
            .O(N__24509),
            .I(N__24496));
    CEMux I__3629 (
            .O(N__24508),
            .I(N__24493));
    CEMux I__3628 (
            .O(N__24507),
            .I(N__24489));
    CEMux I__3627 (
            .O(N__24506),
            .I(N__24486));
    LocalMux I__3626 (
            .O(N__24503),
            .I(N__24480));
    CEMux I__3625 (
            .O(N__24502),
            .I(N__24477));
    CEMux I__3624 (
            .O(N__24501),
            .I(N__24472));
    CEMux I__3623 (
            .O(N__24500),
            .I(N__24469));
    CEMux I__3622 (
            .O(N__24499),
            .I(N__24462));
    LocalMux I__3621 (
            .O(N__24496),
            .I(N__24459));
    LocalMux I__3620 (
            .O(N__24493),
            .I(N__24456));
    CEMux I__3619 (
            .O(N__24492),
            .I(N__24453));
    LocalMux I__3618 (
            .O(N__24489),
            .I(N__24450));
    LocalMux I__3617 (
            .O(N__24486),
            .I(N__24447));
    CEMux I__3616 (
            .O(N__24485),
            .I(N__24444));
    CEMux I__3615 (
            .O(N__24484),
            .I(N__24441));
    CEMux I__3614 (
            .O(N__24483),
            .I(N__24438));
    Span4Mux_s3_h I__3613 (
            .O(N__24480),
            .I(N__24433));
    LocalMux I__3612 (
            .O(N__24477),
            .I(N__24433));
    CEMux I__3611 (
            .O(N__24476),
            .I(N__24430));
    CEMux I__3610 (
            .O(N__24475),
            .I(N__24427));
    LocalMux I__3609 (
            .O(N__24472),
            .I(N__24424));
    LocalMux I__3608 (
            .O(N__24469),
            .I(N__24421));
    CEMux I__3607 (
            .O(N__24468),
            .I(N__24418));
    CEMux I__3606 (
            .O(N__24467),
            .I(N__24415));
    CEMux I__3605 (
            .O(N__24466),
            .I(N__24412));
    CEMux I__3604 (
            .O(N__24465),
            .I(N__24408));
    LocalMux I__3603 (
            .O(N__24462),
            .I(N__24404));
    Span4Mux_v I__3602 (
            .O(N__24459),
            .I(N__24397));
    Span4Mux_v I__3601 (
            .O(N__24456),
            .I(N__24397));
    LocalMux I__3600 (
            .O(N__24453),
            .I(N__24397));
    Span4Mux_h I__3599 (
            .O(N__24450),
            .I(N__24394));
    Span4Mux_h I__3598 (
            .O(N__24447),
            .I(N__24391));
    LocalMux I__3597 (
            .O(N__24444),
            .I(N__24388));
    LocalMux I__3596 (
            .O(N__24441),
            .I(N__24385));
    LocalMux I__3595 (
            .O(N__24438),
            .I(N__24382));
    Span4Mux_h I__3594 (
            .O(N__24433),
            .I(N__24377));
    LocalMux I__3593 (
            .O(N__24430),
            .I(N__24377));
    LocalMux I__3592 (
            .O(N__24427),
            .I(N__24374));
    Span4Mux_h I__3591 (
            .O(N__24424),
            .I(N__24371));
    Span4Mux_s3_h I__3590 (
            .O(N__24421),
            .I(N__24366));
    LocalMux I__3589 (
            .O(N__24418),
            .I(N__24366));
    LocalMux I__3588 (
            .O(N__24415),
            .I(N__24363));
    LocalMux I__3587 (
            .O(N__24412),
            .I(N__24360));
    CEMux I__3586 (
            .O(N__24411),
            .I(N__24357));
    LocalMux I__3585 (
            .O(N__24408),
            .I(N__24354));
    CEMux I__3584 (
            .O(N__24407),
            .I(N__24351));
    Span4Mux_h I__3583 (
            .O(N__24404),
            .I(N__24348));
    Span4Mux_v I__3582 (
            .O(N__24397),
            .I(N__24345));
    Span4Mux_v I__3581 (
            .O(N__24394),
            .I(N__24336));
    Span4Mux_v I__3580 (
            .O(N__24391),
            .I(N__24336));
    Span4Mux_h I__3579 (
            .O(N__24388),
            .I(N__24336));
    Span4Mux_h I__3578 (
            .O(N__24385),
            .I(N__24336));
    Span4Mux_s3_h I__3577 (
            .O(N__24382),
            .I(N__24333));
    Span4Mux_v I__3576 (
            .O(N__24377),
            .I(N__24328));
    Span4Mux_h I__3575 (
            .O(N__24374),
            .I(N__24328));
    Span4Mux_v I__3574 (
            .O(N__24371),
            .I(N__24317));
    Span4Mux_h I__3573 (
            .O(N__24366),
            .I(N__24317));
    Span4Mux_h I__3572 (
            .O(N__24363),
            .I(N__24317));
    Span4Mux_h I__3571 (
            .O(N__24360),
            .I(N__24317));
    LocalMux I__3570 (
            .O(N__24357),
            .I(N__24317));
    Span4Mux_s3_h I__3569 (
            .O(N__24354),
            .I(N__24312));
    LocalMux I__3568 (
            .O(N__24351),
            .I(N__24312));
    Sp12to4 I__3567 (
            .O(N__24348),
            .I(N__24309));
    Span4Mux_v I__3566 (
            .O(N__24345),
            .I(N__24306));
    Span4Mux_v I__3565 (
            .O(N__24336),
            .I(N__24301));
    Span4Mux_h I__3564 (
            .O(N__24333),
            .I(N__24301));
    Span4Mux_v I__3563 (
            .O(N__24328),
            .I(N__24298));
    Span4Mux_v I__3562 (
            .O(N__24317),
            .I(N__24293));
    Span4Mux_h I__3561 (
            .O(N__24312),
            .I(N__24293));
    Odrv12 I__3560 (
            .O(N__24309),
            .I(N_655_g));
    Odrv4 I__3559 (
            .O(N__24306),
            .I(N_655_g));
    Odrv4 I__3558 (
            .O(N__24301),
            .I(N_655_g));
    Odrv4 I__3557 (
            .O(N__24298),
            .I(N_655_g));
    Odrv4 I__3556 (
            .O(N__24293),
            .I(N_655_g));
    InMux I__3555 (
            .O(N__24282),
            .I(N__24278));
    CascadeMux I__3554 (
            .O(N__24281),
            .I(N__24275));
    LocalMux I__3553 (
            .O(N__24278),
            .I(N__24272));
    InMux I__3552 (
            .O(N__24275),
            .I(N__24269));
    Span4Mux_v I__3551 (
            .O(N__24272),
            .I(N__24264));
    LocalMux I__3550 (
            .O(N__24269),
            .I(N__24264));
    Span4Mux_h I__3549 (
            .O(N__24264),
            .I(N__24261));
    Odrv4 I__3548 (
            .O(N__24261),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    CascadeMux I__3547 (
            .O(N__24258),
            .I(N__24254));
    InMux I__3546 (
            .O(N__24257),
            .I(N__24251));
    InMux I__3545 (
            .O(N__24254),
            .I(N__24248));
    LocalMux I__3544 (
            .O(N__24251),
            .I(N__24243));
    LocalMux I__3543 (
            .O(N__24248),
            .I(N__24243));
    Span4Mux_h I__3542 (
            .O(N__24243),
            .I(N__24240));
    Odrv4 I__3541 (
            .O(N__24240),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    InMux I__3540 (
            .O(N__24237),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    InMux I__3539 (
            .O(N__24234),
            .I(N__24230));
    CascadeMux I__3538 (
            .O(N__24233),
            .I(N__24227));
    LocalMux I__3537 (
            .O(N__24230),
            .I(N__24224));
    InMux I__3536 (
            .O(N__24227),
            .I(N__24221));
    Span4Mux_v I__3535 (
            .O(N__24224),
            .I(N__24216));
    LocalMux I__3534 (
            .O(N__24221),
            .I(N__24216));
    Span4Mux_h I__3533 (
            .O(N__24216),
            .I(N__24213));
    Odrv4 I__3532 (
            .O(N__24213),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__3531 (
            .O(N__24210),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    CascadeMux I__3530 (
            .O(N__24207),
            .I(N__24203));
    InMux I__3529 (
            .O(N__24206),
            .I(N__24200));
    InMux I__3528 (
            .O(N__24203),
            .I(N__24197));
    LocalMux I__3527 (
            .O(N__24200),
            .I(N__24194));
    LocalMux I__3526 (
            .O(N__24197),
            .I(N__24191));
    Span4Mux_v I__3525 (
            .O(N__24194),
            .I(N__24186));
    Span4Mux_v I__3524 (
            .O(N__24191),
            .I(N__24186));
    Odrv4 I__3523 (
            .O(N__24186),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__3522 (
            .O(N__24183),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    InMux I__3521 (
            .O(N__24180),
            .I(N__24175));
    InMux I__3520 (
            .O(N__24179),
            .I(N__24172));
    InMux I__3519 (
            .O(N__24178),
            .I(N__24169));
    LocalMux I__3518 (
            .O(N__24175),
            .I(N__24166));
    LocalMux I__3517 (
            .O(N__24172),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__3516 (
            .O(N__24169),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__3515 (
            .O(N__24166),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__3514 (
            .O(N__24159),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__3513 (
            .O(N__24156),
            .I(N__24151));
    InMux I__3512 (
            .O(N__24155),
            .I(N__24148));
    InMux I__3511 (
            .O(N__24154),
            .I(N__24145));
    LocalMux I__3510 (
            .O(N__24151),
            .I(N__24142));
    LocalMux I__3509 (
            .O(N__24148),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__3508 (
            .O(N__24145),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__3507 (
            .O(N__24142),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__3506 (
            .O(N__24135),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__3505 (
            .O(N__24132),
            .I(N__24127));
    InMux I__3504 (
            .O(N__24131),
            .I(N__24124));
    InMux I__3503 (
            .O(N__24130),
            .I(N__24121));
    LocalMux I__3502 (
            .O(N__24127),
            .I(N__24118));
    LocalMux I__3501 (
            .O(N__24124),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__3500 (
            .O(N__24121),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__3499 (
            .O(N__24118),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__3498 (
            .O(N__24111),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__3497 (
            .O(N__24108),
            .I(N__24103));
    InMux I__3496 (
            .O(N__24107),
            .I(N__24100));
    InMux I__3495 (
            .O(N__24106),
            .I(N__24097));
    LocalMux I__3494 (
            .O(N__24103),
            .I(N__24094));
    LocalMux I__3493 (
            .O(N__24100),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__3492 (
            .O(N__24097),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__3491 (
            .O(N__24094),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__3490 (
            .O(N__24087),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__3489 (
            .O(N__24084),
            .I(N__24080));
    InMux I__3488 (
            .O(N__24083),
            .I(N__24076));
    LocalMux I__3487 (
            .O(N__24080),
            .I(N__24073));
    InMux I__3486 (
            .O(N__24079),
            .I(N__24070));
    LocalMux I__3485 (
            .O(N__24076),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__3484 (
            .O(N__24073),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__3483 (
            .O(N__24070),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__3482 (
            .O(N__24063),
            .I(bfn_8_9_0_));
    InMux I__3481 (
            .O(N__24060),
            .I(N__24048));
    InMux I__3480 (
            .O(N__24059),
            .I(N__24048));
    InMux I__3479 (
            .O(N__24058),
            .I(N__24048));
    InMux I__3478 (
            .O(N__24057),
            .I(N__24048));
    LocalMux I__3477 (
            .O(N__24048),
            .I(N__24039));
    InMux I__3476 (
            .O(N__24047),
            .I(N__24034));
    InMux I__3475 (
            .O(N__24046),
            .I(N__24034));
    InMux I__3474 (
            .O(N__24045),
            .I(N__24025));
    InMux I__3473 (
            .O(N__24044),
            .I(N__24025));
    InMux I__3472 (
            .O(N__24043),
            .I(N__24025));
    InMux I__3471 (
            .O(N__24042),
            .I(N__24025));
    Odrv4 I__3470 (
            .O(N__24039),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__3469 (
            .O(N__24034),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__3468 (
            .O(N__24025),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__3467 (
            .O(N__24018),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__3466 (
            .O(N__24015),
            .I(N__24011));
    InMux I__3465 (
            .O(N__24014),
            .I(N__24007));
    LocalMux I__3464 (
            .O(N__24011),
            .I(N__24004));
    InMux I__3463 (
            .O(N__24010),
            .I(N__24001));
    LocalMux I__3462 (
            .O(N__24007),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__3461 (
            .O(N__24004),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__3460 (
            .O(N__24001),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__3459 (
            .O(N__23994),
            .I(N__23990));
    InMux I__3458 (
            .O(N__23993),
            .I(N__23987));
    LocalMux I__3457 (
            .O(N__23990),
            .I(N__23984));
    LocalMux I__3456 (
            .O(N__23987),
            .I(N__23981));
    Odrv4 I__3455 (
            .O(N__23984),
            .I(\current_shift_inst.PI_CTRL.N_47_16 ));
    Odrv4 I__3454 (
            .O(N__23981),
            .I(\current_shift_inst.PI_CTRL.N_47_16 ));
    InMux I__3453 (
            .O(N__23976),
            .I(N__23972));
    InMux I__3452 (
            .O(N__23975),
            .I(N__23969));
    LocalMux I__3451 (
            .O(N__23972),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    LocalMux I__3450 (
            .O(N__23969),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    InMux I__3449 (
            .O(N__23964),
            .I(N__23958));
    CascadeMux I__3448 (
            .O(N__23963),
            .I(N__23955));
    CascadeMux I__3447 (
            .O(N__23962),
            .I(N__23952));
    InMux I__3446 (
            .O(N__23961),
            .I(N__23948));
    LocalMux I__3445 (
            .O(N__23958),
            .I(N__23945));
    InMux I__3444 (
            .O(N__23955),
            .I(N__23941));
    InMux I__3443 (
            .O(N__23952),
            .I(N__23936));
    InMux I__3442 (
            .O(N__23951),
            .I(N__23936));
    LocalMux I__3441 (
            .O(N__23948),
            .I(N__23933));
    Span4Mux_v I__3440 (
            .O(N__23945),
            .I(N__23930));
    InMux I__3439 (
            .O(N__23944),
            .I(N__23927));
    LocalMux I__3438 (
            .O(N__23941),
            .I(N__23922));
    LocalMux I__3437 (
            .O(N__23936),
            .I(N__23922));
    Span4Mux_h I__3436 (
            .O(N__23933),
            .I(N__23915));
    Span4Mux_h I__3435 (
            .O(N__23930),
            .I(N__23915));
    LocalMux I__3434 (
            .O(N__23927),
            .I(N__23915));
    Span4Mux_h I__3433 (
            .O(N__23922),
            .I(N__23912));
    Span4Mux_v I__3432 (
            .O(N__23915),
            .I(N__23909));
    Odrv4 I__3431 (
            .O(N__23912),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__3430 (
            .O(N__23909),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__3429 (
            .O(N__23904),
            .I(N__23899));
    InMux I__3428 (
            .O(N__23903),
            .I(N__23895));
    InMux I__3427 (
            .O(N__23902),
            .I(N__23892));
    InMux I__3426 (
            .O(N__23899),
            .I(N__23889));
    CascadeMux I__3425 (
            .O(N__23898),
            .I(N__23886));
    LocalMux I__3424 (
            .O(N__23895),
            .I(N__23883));
    LocalMux I__3423 (
            .O(N__23892),
            .I(N__23880));
    LocalMux I__3422 (
            .O(N__23889),
            .I(N__23877));
    InMux I__3421 (
            .O(N__23886),
            .I(N__23874));
    Span12Mux_v I__3420 (
            .O(N__23883),
            .I(N__23871));
    Span4Mux_v I__3419 (
            .O(N__23880),
            .I(N__23868));
    Odrv4 I__3418 (
            .O(N__23877),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__3417 (
            .O(N__23874),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv12 I__3416 (
            .O(N__23871),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__3415 (
            .O(N__23868),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__3414 (
            .O(N__23859),
            .I(N__23856));
    LocalMux I__3413 (
            .O(N__23856),
            .I(N__23850));
    InMux I__3412 (
            .O(N__23855),
            .I(N__23847));
    InMux I__3411 (
            .O(N__23854),
            .I(N__23844));
    InMux I__3410 (
            .O(N__23853),
            .I(N__23841));
    Span4Mux_v I__3409 (
            .O(N__23850),
            .I(N__23836));
    LocalMux I__3408 (
            .O(N__23847),
            .I(N__23836));
    LocalMux I__3407 (
            .O(N__23844),
            .I(N__23833));
    LocalMux I__3406 (
            .O(N__23841),
            .I(N__23830));
    Odrv4 I__3405 (
            .O(N__23836),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__3404 (
            .O(N__23833),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__3403 (
            .O(N__23830),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__3402 (
            .O(N__23823),
            .I(N__23819));
    InMux I__3401 (
            .O(N__23822),
            .I(N__23815));
    InMux I__3400 (
            .O(N__23819),
            .I(N__23812));
    InMux I__3399 (
            .O(N__23818),
            .I(N__23809));
    LocalMux I__3398 (
            .O(N__23815),
            .I(N__23805));
    LocalMux I__3397 (
            .O(N__23812),
            .I(N__23800));
    LocalMux I__3396 (
            .O(N__23809),
            .I(N__23800));
    InMux I__3395 (
            .O(N__23808),
            .I(N__23797));
    Span4Mux_v I__3394 (
            .O(N__23805),
            .I(N__23792));
    Span4Mux_v I__3393 (
            .O(N__23800),
            .I(N__23792));
    LocalMux I__3392 (
            .O(N__23797),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__3391 (
            .O(N__23792),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    CascadeMux I__3390 (
            .O(N__23787),
            .I(N__23784));
    InMux I__3389 (
            .O(N__23784),
            .I(N__23780));
    CascadeMux I__3388 (
            .O(N__23783),
            .I(N__23776));
    LocalMux I__3387 (
            .O(N__23780),
            .I(N__23772));
    InMux I__3386 (
            .O(N__23779),
            .I(N__23769));
    InMux I__3385 (
            .O(N__23776),
            .I(N__23766));
    InMux I__3384 (
            .O(N__23775),
            .I(N__23763));
    Span4Mux_v I__3383 (
            .O(N__23772),
            .I(N__23758));
    LocalMux I__3382 (
            .O(N__23769),
            .I(N__23758));
    LocalMux I__3381 (
            .O(N__23766),
            .I(N__23755));
    LocalMux I__3380 (
            .O(N__23763),
            .I(N__23752));
    Odrv4 I__3379 (
            .O(N__23758),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__3378 (
            .O(N__23755),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__3377 (
            .O(N__23752),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__3376 (
            .O(N__23745),
            .I(N__23742));
    LocalMux I__3375 (
            .O(N__23742),
            .I(N__23739));
    Span4Mux_v I__3374 (
            .O(N__23739),
            .I(N__23736));
    Odrv4 I__3373 (
            .O(N__23736),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    CascadeMux I__3372 (
            .O(N__23733),
            .I(N__23730));
    InMux I__3371 (
            .O(N__23730),
            .I(N__23727));
    LocalMux I__3370 (
            .O(N__23727),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__3369 (
            .O(N__23724),
            .I(N__23721));
    InMux I__3368 (
            .O(N__23721),
            .I(N__23718));
    LocalMux I__3367 (
            .O(N__23718),
            .I(N__23715));
    Odrv4 I__3366 (
            .O(N__23715),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__3365 (
            .O(N__23712),
            .I(N__23709));
    LocalMux I__3364 (
            .O(N__23709),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__3363 (
            .O(N__23706),
            .I(N__23703));
    InMux I__3362 (
            .O(N__23703),
            .I(N__23700));
    LocalMux I__3361 (
            .O(N__23700),
            .I(N__23697));
    Span4Mux_v I__3360 (
            .O(N__23697),
            .I(N__23694));
    Odrv4 I__3359 (
            .O(N__23694),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__3358 (
            .O(N__23691),
            .I(N__23688));
    LocalMux I__3357 (
            .O(N__23688),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__3356 (
            .O(N__23685),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__3355 (
            .O(N__23682),
            .I(N__23679));
    LocalMux I__3354 (
            .O(N__23679),
            .I(N__23676));
    IoSpan4Mux I__3353 (
            .O(N__23676),
            .I(N__23673));
    Span4Mux_s2_v I__3352 (
            .O(N__23673),
            .I(N__23670));
    Span4Mux_v I__3351 (
            .O(N__23670),
            .I(N__23667));
    Span4Mux_h I__3350 (
            .O(N__23667),
            .I(N__23664));
    Span4Mux_h I__3349 (
            .O(N__23664),
            .I(N__23661));
    Odrv4 I__3348 (
            .O(N__23661),
            .I(pwm_output_c));
    InMux I__3347 (
            .O(N__23658),
            .I(N__23654));
    InMux I__3346 (
            .O(N__23657),
            .I(N__23650));
    LocalMux I__3345 (
            .O(N__23654),
            .I(N__23647));
    InMux I__3344 (
            .O(N__23653),
            .I(N__23644));
    LocalMux I__3343 (
            .O(N__23650),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__3342 (
            .O(N__23647),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__3341 (
            .O(N__23644),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__3340 (
            .O(N__23637),
            .I(bfn_8_8_0_));
    InMux I__3339 (
            .O(N__23634),
            .I(N__23629));
    InMux I__3338 (
            .O(N__23633),
            .I(N__23626));
    InMux I__3337 (
            .O(N__23632),
            .I(N__23623));
    LocalMux I__3336 (
            .O(N__23629),
            .I(N__23620));
    LocalMux I__3335 (
            .O(N__23626),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__3334 (
            .O(N__23623),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__3333 (
            .O(N__23620),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__3332 (
            .O(N__23613),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__3331 (
            .O(N__23610),
            .I(N__23606));
    InMux I__3330 (
            .O(N__23609),
            .I(N__23602));
    LocalMux I__3329 (
            .O(N__23606),
            .I(N__23599));
    InMux I__3328 (
            .O(N__23605),
            .I(N__23596));
    LocalMux I__3327 (
            .O(N__23602),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__3326 (
            .O(N__23599),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__3325 (
            .O(N__23596),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__3324 (
            .O(N__23589),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__3323 (
            .O(N__23586),
            .I(N__23581));
    InMux I__3322 (
            .O(N__23585),
            .I(N__23578));
    InMux I__3321 (
            .O(N__23584),
            .I(N__23575));
    LocalMux I__3320 (
            .O(N__23581),
            .I(N__23572));
    LocalMux I__3319 (
            .O(N__23578),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__3318 (
            .O(N__23575),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__3317 (
            .O(N__23572),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__3316 (
            .O(N__23565),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__3315 (
            .O(N__23562),
            .I(N__23559));
    LocalMux I__3314 (
            .O(N__23559),
            .I(N__23556));
    Odrv12 I__3313 (
            .O(N__23556),
            .I(il_max_comp1_c));
    CascadeMux I__3312 (
            .O(N__23553),
            .I(N__23550));
    InMux I__3311 (
            .O(N__23550),
            .I(N__23547));
    LocalMux I__3310 (
            .O(N__23547),
            .I(N__23544));
    Span4Mux_v I__3309 (
            .O(N__23544),
            .I(N__23541));
    Span4Mux_h I__3308 (
            .O(N__23541),
            .I(N__23538));
    Odrv4 I__3307 (
            .O(N__23538),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    InMux I__3306 (
            .O(N__23535),
            .I(N__23532));
    LocalMux I__3305 (
            .O(N__23532),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__3304 (
            .O(N__23529),
            .I(N__23526));
    InMux I__3303 (
            .O(N__23526),
            .I(N__23523));
    LocalMux I__3302 (
            .O(N__23523),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    InMux I__3301 (
            .O(N__23520),
            .I(N__23517));
    LocalMux I__3300 (
            .O(N__23517),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__3299 (
            .O(N__23514),
            .I(N__23511));
    InMux I__3298 (
            .O(N__23511),
            .I(N__23508));
    LocalMux I__3297 (
            .O(N__23508),
            .I(N__23505));
    Odrv4 I__3296 (
            .O(N__23505),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    InMux I__3295 (
            .O(N__23502),
            .I(N__23499));
    LocalMux I__3294 (
            .O(N__23499),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__3293 (
            .O(N__23496),
            .I(N__23493));
    LocalMux I__3292 (
            .O(N__23493),
            .I(N__23490));
    Span4Mux_h I__3291 (
            .O(N__23490),
            .I(N__23487));
    Odrv4 I__3290 (
            .O(N__23487),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    CascadeMux I__3289 (
            .O(N__23484),
            .I(N__23481));
    InMux I__3288 (
            .O(N__23481),
            .I(N__23478));
    LocalMux I__3287 (
            .O(N__23478),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__3286 (
            .O(N__23475),
            .I(N__23472));
    InMux I__3285 (
            .O(N__23472),
            .I(N__23469));
    LocalMux I__3284 (
            .O(N__23469),
            .I(N__23466));
    Odrv4 I__3283 (
            .O(N__23466),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    InMux I__3282 (
            .O(N__23463),
            .I(N__23460));
    LocalMux I__3281 (
            .O(N__23460),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__3280 (
            .O(N__23457),
            .I(N__23454));
    InMux I__3279 (
            .O(N__23454),
            .I(N__23451));
    LocalMux I__3278 (
            .O(N__23451),
            .I(N__23448));
    Span4Mux_v I__3277 (
            .O(N__23448),
            .I(N__23445));
    Odrv4 I__3276 (
            .O(N__23445),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    InMux I__3275 (
            .O(N__23442),
            .I(N__23439));
    LocalMux I__3274 (
            .O(N__23439),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__3273 (
            .O(N__23436),
            .I(N__23433));
    InMux I__3272 (
            .O(N__23433),
            .I(N__23430));
    LocalMux I__3271 (
            .O(N__23430),
            .I(N__23427));
    Odrv12 I__3270 (
            .O(N__23427),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__3269 (
            .O(N__23424),
            .I(N__23421));
    LocalMux I__3268 (
            .O(N__23421),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__3267 (
            .O(N__23418),
            .I(\current_shift_inst.timer_phase.counter_cry_20 ));
    InMux I__3266 (
            .O(N__23415),
            .I(\current_shift_inst.timer_phase.counter_cry_21 ));
    InMux I__3265 (
            .O(N__23412),
            .I(\current_shift_inst.timer_phase.counter_cry_22 ));
    InMux I__3264 (
            .O(N__23409),
            .I(bfn_7_22_0_));
    InMux I__3263 (
            .O(N__23406),
            .I(\current_shift_inst.timer_phase.counter_cry_24 ));
    InMux I__3262 (
            .O(N__23403),
            .I(\current_shift_inst.timer_phase.counter_cry_25 ));
    InMux I__3261 (
            .O(N__23400),
            .I(\current_shift_inst.timer_phase.counter_cry_26 ));
    InMux I__3260 (
            .O(N__23397),
            .I(\current_shift_inst.timer_phase.counter_cry_27 ));
    InMux I__3259 (
            .O(N__23394),
            .I(\current_shift_inst.timer_phase.counter_cry_28 ));
    InMux I__3258 (
            .O(N__23391),
            .I(N__23388));
    LocalMux I__3257 (
            .O(N__23388),
            .I(N__23385));
    Span4Mux_h I__3256 (
            .O(N__23385),
            .I(N__23382));
    Odrv4 I__3255 (
            .O(N__23382),
            .I(il_min_comp2_c));
    InMux I__3254 (
            .O(N__23379),
            .I(\current_shift_inst.timer_phase.counter_cry_11 ));
    InMux I__3253 (
            .O(N__23376),
            .I(\current_shift_inst.timer_phase.counter_cry_12 ));
    InMux I__3252 (
            .O(N__23373),
            .I(\current_shift_inst.timer_phase.counter_cry_13 ));
    InMux I__3251 (
            .O(N__23370),
            .I(\current_shift_inst.timer_phase.counter_cry_14 ));
    InMux I__3250 (
            .O(N__23367),
            .I(bfn_7_21_0_));
    InMux I__3249 (
            .O(N__23364),
            .I(\current_shift_inst.timer_phase.counter_cry_16 ));
    InMux I__3248 (
            .O(N__23361),
            .I(\current_shift_inst.timer_phase.counter_cry_17 ));
    InMux I__3247 (
            .O(N__23358),
            .I(\current_shift_inst.timer_phase.counter_cry_18 ));
    InMux I__3246 (
            .O(N__23355),
            .I(\current_shift_inst.timer_phase.counter_cry_19 ));
    InMux I__3245 (
            .O(N__23352),
            .I(\current_shift_inst.timer_phase.counter_cry_2 ));
    InMux I__3244 (
            .O(N__23349),
            .I(\current_shift_inst.timer_phase.counter_cry_3 ));
    InMux I__3243 (
            .O(N__23346),
            .I(\current_shift_inst.timer_phase.counter_cry_4 ));
    InMux I__3242 (
            .O(N__23343),
            .I(\current_shift_inst.timer_phase.counter_cry_5 ));
    InMux I__3241 (
            .O(N__23340),
            .I(\current_shift_inst.timer_phase.counter_cry_6 ));
    InMux I__3240 (
            .O(N__23337),
            .I(bfn_7_20_0_));
    InMux I__3239 (
            .O(N__23334),
            .I(\current_shift_inst.timer_phase.counter_cry_8 ));
    InMux I__3238 (
            .O(N__23331),
            .I(\current_shift_inst.timer_phase.counter_cry_9 ));
    InMux I__3237 (
            .O(N__23328),
            .I(\current_shift_inst.timer_phase.counter_cry_10 ));
    InMux I__3236 (
            .O(N__23325),
            .I(bfn_7_19_0_));
    InMux I__3235 (
            .O(N__23322),
            .I(\current_shift_inst.timer_phase.counter_cry_0 ));
    InMux I__3234 (
            .O(N__23319),
            .I(\current_shift_inst.timer_phase.counter_cry_1 ));
    CascadeMux I__3233 (
            .O(N__23316),
            .I(N__23313));
    InMux I__3232 (
            .O(N__23313),
            .I(N__23310));
    LocalMux I__3231 (
            .O(N__23310),
            .I(N__23307));
    Sp12to4 I__3230 (
            .O(N__23307),
            .I(N__23304));
    Odrv12 I__3229 (
            .O(N__23304),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__3228 (
            .O(N__23301),
            .I(N__23298));
    LocalMux I__3227 (
            .O(N__23298),
            .I(N__23295));
    Odrv12 I__3226 (
            .O(N__23295),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__3225 (
            .O(N__23292),
            .I(N__23289));
    LocalMux I__3224 (
            .O(N__23289),
            .I(N__23284));
    InMux I__3223 (
            .O(N__23288),
            .I(N__23281));
    CascadeMux I__3222 (
            .O(N__23287),
            .I(N__23277));
    Span4Mux_v I__3221 (
            .O(N__23284),
            .I(N__23272));
    LocalMux I__3220 (
            .O(N__23281),
            .I(N__23272));
    InMux I__3219 (
            .O(N__23280),
            .I(N__23267));
    InMux I__3218 (
            .O(N__23277),
            .I(N__23267));
    Odrv4 I__3217 (
            .O(N__23272),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__3216 (
            .O(N__23267),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__3215 (
            .O(N__23262),
            .I(N__23259));
    LocalMux I__3214 (
            .O(N__23259),
            .I(N__23254));
    InMux I__3213 (
            .O(N__23258),
            .I(N__23251));
    InMux I__3212 (
            .O(N__23257),
            .I(N__23247));
    Span4Mux_v I__3211 (
            .O(N__23254),
            .I(N__23242));
    LocalMux I__3210 (
            .O(N__23251),
            .I(N__23242));
    InMux I__3209 (
            .O(N__23250),
            .I(N__23239));
    LocalMux I__3208 (
            .O(N__23247),
            .I(N__23236));
    Span4Mux_v I__3207 (
            .O(N__23242),
            .I(N__23233));
    LocalMux I__3206 (
            .O(N__23239),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv12 I__3205 (
            .O(N__23236),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__3204 (
            .O(N__23233),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__3203 (
            .O(N__23226),
            .I(N__23221));
    InMux I__3202 (
            .O(N__23225),
            .I(N__23217));
    InMux I__3201 (
            .O(N__23224),
            .I(N__23214));
    LocalMux I__3200 (
            .O(N__23221),
            .I(N__23211));
    InMux I__3199 (
            .O(N__23220),
            .I(N__23208));
    LocalMux I__3198 (
            .O(N__23217),
            .I(N__23205));
    LocalMux I__3197 (
            .O(N__23214),
            .I(N__23202));
    Span4Mux_v I__3196 (
            .O(N__23211),
            .I(N__23195));
    LocalMux I__3195 (
            .O(N__23208),
            .I(N__23195));
    Span4Mux_h I__3194 (
            .O(N__23205),
            .I(N__23195));
    Odrv4 I__3193 (
            .O(N__23202),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__3192 (
            .O(N__23195),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__3191 (
            .O(N__23190),
            .I(N__23185));
    CascadeMux I__3190 (
            .O(N__23189),
            .I(N__23182));
    CascadeMux I__3189 (
            .O(N__23188),
            .I(N__23179));
    InMux I__3188 (
            .O(N__23185),
            .I(N__23176));
    InMux I__3187 (
            .O(N__23182),
            .I(N__23172));
    InMux I__3186 (
            .O(N__23179),
            .I(N__23169));
    LocalMux I__3185 (
            .O(N__23176),
            .I(N__23166));
    InMux I__3184 (
            .O(N__23175),
            .I(N__23163));
    LocalMux I__3183 (
            .O(N__23172),
            .I(N__23160));
    LocalMux I__3182 (
            .O(N__23169),
            .I(N__23157));
    Span4Mux_v I__3181 (
            .O(N__23166),
            .I(N__23150));
    LocalMux I__3180 (
            .O(N__23163),
            .I(N__23150));
    Span4Mux_h I__3179 (
            .O(N__23160),
            .I(N__23150));
    Odrv4 I__3178 (
            .O(N__23157),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__3177 (
            .O(N__23150),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__3176 (
            .O(N__23145),
            .I(N__23139));
    CascadeMux I__3175 (
            .O(N__23144),
            .I(N__23136));
    InMux I__3174 (
            .O(N__23143),
            .I(N__23133));
    InMux I__3173 (
            .O(N__23142),
            .I(N__23130));
    LocalMux I__3172 (
            .O(N__23139),
            .I(N__23127));
    InMux I__3171 (
            .O(N__23136),
            .I(N__23124));
    LocalMux I__3170 (
            .O(N__23133),
            .I(N__23121));
    LocalMux I__3169 (
            .O(N__23130),
            .I(N__23118));
    Span4Mux_v I__3168 (
            .O(N__23127),
            .I(N__23111));
    LocalMux I__3167 (
            .O(N__23124),
            .I(N__23111));
    Span4Mux_h I__3166 (
            .O(N__23121),
            .I(N__23111));
    Odrv4 I__3165 (
            .O(N__23118),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__3164 (
            .O(N__23111),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__3163 (
            .O(N__23106),
            .I(N__23101));
    InMux I__3162 (
            .O(N__23105),
            .I(N__23095));
    InMux I__3161 (
            .O(N__23104),
            .I(N__23095));
    LocalMux I__3160 (
            .O(N__23101),
            .I(N__23092));
    InMux I__3159 (
            .O(N__23100),
            .I(N__23089));
    LocalMux I__3158 (
            .O(N__23095),
            .I(N__23086));
    Odrv12 I__3157 (
            .O(N__23092),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__3156 (
            .O(N__23089),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__3155 (
            .O(N__23086),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__3154 (
            .O(N__23079),
            .I(N__23076));
    InMux I__3153 (
            .O(N__23076),
            .I(N__23068));
    InMux I__3152 (
            .O(N__23075),
            .I(N__23068));
    InMux I__3151 (
            .O(N__23074),
            .I(N__23065));
    InMux I__3150 (
            .O(N__23073),
            .I(N__23062));
    LocalMux I__3149 (
            .O(N__23068),
            .I(N__23059));
    LocalMux I__3148 (
            .O(N__23065),
            .I(N__23056));
    LocalMux I__3147 (
            .O(N__23062),
            .I(N__23051));
    Span4Mux_h I__3146 (
            .O(N__23059),
            .I(N__23051));
    Odrv12 I__3145 (
            .O(N__23056),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__3144 (
            .O(N__23051),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__3143 (
            .O(N__23046),
            .I(N__23041));
    InMux I__3142 (
            .O(N__23045),
            .I(N__23038));
    InMux I__3141 (
            .O(N__23044),
            .I(N__23032));
    InMux I__3140 (
            .O(N__23041),
            .I(N__23032));
    LocalMux I__3139 (
            .O(N__23038),
            .I(N__23029));
    InMux I__3138 (
            .O(N__23037),
            .I(N__23026));
    LocalMux I__3137 (
            .O(N__23032),
            .I(N__23023));
    Odrv4 I__3136 (
            .O(N__23029),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__3135 (
            .O(N__23026),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__3134 (
            .O(N__23023),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__3133 (
            .O(N__23016),
            .I(N__23012));
    InMux I__3132 (
            .O(N__23015),
            .I(N__23009));
    LocalMux I__3131 (
            .O(N__23012),
            .I(N__23006));
    LocalMux I__3130 (
            .O(N__23009),
            .I(N__23003));
    Odrv12 I__3129 (
            .O(N__23006),
            .I(\current_shift_inst.PI_CTRL.N_46_16 ));
    Odrv4 I__3128 (
            .O(N__23003),
            .I(\current_shift_inst.PI_CTRL.N_46_16 ));
    CascadeMux I__3127 (
            .O(N__22998),
            .I(N__22995));
    InMux I__3126 (
            .O(N__22995),
            .I(N__22992));
    LocalMux I__3125 (
            .O(N__22992),
            .I(N__22989));
    Span4Mux_h I__3124 (
            .O(N__22989),
            .I(N__22986));
    Odrv4 I__3123 (
            .O(N__22986),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__3122 (
            .O(N__22983),
            .I(N__22979));
    CascadeMux I__3121 (
            .O(N__22982),
            .I(N__22975));
    LocalMux I__3120 (
            .O(N__22979),
            .I(N__22971));
    InMux I__3119 (
            .O(N__22978),
            .I(N__22968));
    InMux I__3118 (
            .O(N__22975),
            .I(N__22965));
    CascadeMux I__3117 (
            .O(N__22974),
            .I(N__22962));
    Span4Mux_v I__3116 (
            .O(N__22971),
            .I(N__22957));
    LocalMux I__3115 (
            .O(N__22968),
            .I(N__22957));
    LocalMux I__3114 (
            .O(N__22965),
            .I(N__22954));
    InMux I__3113 (
            .O(N__22962),
            .I(N__22951));
    Odrv4 I__3112 (
            .O(N__22957),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__3111 (
            .O(N__22954),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__3110 (
            .O(N__22951),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__3109 (
            .O(N__22944),
            .I(N__22941));
    LocalMux I__3108 (
            .O(N__22941),
            .I(N__22938));
    Odrv12 I__3107 (
            .O(N__22938),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    CascadeMux I__3106 (
            .O(N__22935),
            .I(N__22929));
    CascadeMux I__3105 (
            .O(N__22934),
            .I(N__22926));
    CascadeMux I__3104 (
            .O(N__22933),
            .I(N__22921));
    CascadeMux I__3103 (
            .O(N__22932),
            .I(N__22918));
    InMux I__3102 (
            .O(N__22929),
            .I(N__22910));
    InMux I__3101 (
            .O(N__22926),
            .I(N__22910));
    InMux I__3100 (
            .O(N__22925),
            .I(N__22910));
    InMux I__3099 (
            .O(N__22924),
            .I(N__22901));
    InMux I__3098 (
            .O(N__22921),
            .I(N__22901));
    InMux I__3097 (
            .O(N__22918),
            .I(N__22901));
    InMux I__3096 (
            .O(N__22917),
            .I(N__22901));
    LocalMux I__3095 (
            .O(N__22910),
            .I(N__22896));
    LocalMux I__3094 (
            .O(N__22901),
            .I(N__22896));
    Span4Mux_h I__3093 (
            .O(N__22896),
            .I(N__22893));
    Odrv4 I__3092 (
            .O(N__22893),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    InMux I__3091 (
            .O(N__22890),
            .I(N__22887));
    LocalMux I__3090 (
            .O(N__22887),
            .I(N__22884));
    Odrv4 I__3089 (
            .O(N__22884),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    CascadeMux I__3088 (
            .O(N__22881),
            .I(N__22878));
    InMux I__3087 (
            .O(N__22878),
            .I(N__22875));
    LocalMux I__3086 (
            .O(N__22875),
            .I(N__22872));
    Span4Mux_h I__3085 (
            .O(N__22872),
            .I(N__22869));
    Odrv4 I__3084 (
            .O(N__22869),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    InMux I__3083 (
            .O(N__22866),
            .I(N__22863));
    LocalMux I__3082 (
            .O(N__22863),
            .I(N__22860));
    Odrv4 I__3081 (
            .O(N__22860),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    CascadeMux I__3080 (
            .O(N__22857),
            .I(N__22853));
    InMux I__3079 (
            .O(N__22856),
            .I(N__22850));
    InMux I__3078 (
            .O(N__22853),
            .I(N__22847));
    LocalMux I__3077 (
            .O(N__22850),
            .I(N__22843));
    LocalMux I__3076 (
            .O(N__22847),
            .I(N__22839));
    InMux I__3075 (
            .O(N__22846),
            .I(N__22836));
    Span4Mux_h I__3074 (
            .O(N__22843),
            .I(N__22833));
    InMux I__3073 (
            .O(N__22842),
            .I(N__22830));
    Span4Mux_h I__3072 (
            .O(N__22839),
            .I(N__22825));
    LocalMux I__3071 (
            .O(N__22836),
            .I(N__22825));
    Odrv4 I__3070 (
            .O(N__22833),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__3069 (
            .O(N__22830),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__3068 (
            .O(N__22825),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__3067 (
            .O(N__22818),
            .I(N__22815));
    LocalMux I__3066 (
            .O(N__22815),
            .I(\current_shift_inst.PI_CTRL.N_46_21 ));
    InMux I__3065 (
            .O(N__22812),
            .I(N__22809));
    LocalMux I__3064 (
            .O(N__22809),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_2 ));
    CascadeMux I__3063 (
            .O(N__22806),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2_cascade_ ));
    InMux I__3062 (
            .O(N__22803),
            .I(N__22797));
    InMux I__3061 (
            .O(N__22802),
            .I(N__22790));
    InMux I__3060 (
            .O(N__22801),
            .I(N__22790));
    InMux I__3059 (
            .O(N__22800),
            .I(N__22790));
    LocalMux I__3058 (
            .O(N__22797),
            .I(N__22787));
    LocalMux I__3057 (
            .O(N__22790),
            .I(N__22784));
    Odrv12 I__3056 (
            .O(N__22787),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__3055 (
            .O(N__22784),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    InMux I__3054 (
            .O(N__22779),
            .I(N__22776));
    LocalMux I__3053 (
            .O(N__22776),
            .I(N__22773));
    Odrv4 I__3052 (
            .O(N__22773),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ));
    CascadeMux I__3051 (
            .O(N__22770),
            .I(N__22767));
    InMux I__3050 (
            .O(N__22767),
            .I(N__22764));
    LocalMux I__3049 (
            .O(N__22764),
            .I(N__22761));
    Odrv4 I__3048 (
            .O(N__22761),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ));
    InMux I__3047 (
            .O(N__22758),
            .I(N__22755));
    LocalMux I__3046 (
            .O(N__22755),
            .I(N__22752));
    Odrv12 I__3045 (
            .O(N__22752),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__3044 (
            .O(N__22749),
            .I(N__22746));
    LocalMux I__3043 (
            .O(N__22746),
            .I(N__22743));
    Span4Mux_h I__3042 (
            .O(N__22743),
            .I(N__22740));
    Odrv4 I__3041 (
            .O(N__22740),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__3040 (
            .O(N__22737),
            .I(N__22731));
    InMux I__3039 (
            .O(N__22736),
            .I(N__22728));
    InMux I__3038 (
            .O(N__22735),
            .I(N__22725));
    InMux I__3037 (
            .O(N__22734),
            .I(N__22722));
    LocalMux I__3036 (
            .O(N__22731),
            .I(N__22719));
    LocalMux I__3035 (
            .O(N__22728),
            .I(N__22716));
    LocalMux I__3034 (
            .O(N__22725),
            .I(N__22713));
    LocalMux I__3033 (
            .O(N__22722),
            .I(N__22710));
    Span12Mux_v I__3032 (
            .O(N__22719),
            .I(N__22707));
    Odrv12 I__3031 (
            .O(N__22716),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__3030 (
            .O(N__22713),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__3029 (
            .O(N__22710),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv12 I__3028 (
            .O(N__22707),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__3027 (
            .O(N__22698),
            .I(N__22692));
    InMux I__3026 (
            .O(N__22697),
            .I(N__22689));
    CascadeMux I__3025 (
            .O(N__22696),
            .I(N__22686));
    InMux I__3024 (
            .O(N__22695),
            .I(N__22683));
    LocalMux I__3023 (
            .O(N__22692),
            .I(N__22680));
    LocalMux I__3022 (
            .O(N__22689),
            .I(N__22677));
    InMux I__3021 (
            .O(N__22686),
            .I(N__22674));
    LocalMux I__3020 (
            .O(N__22683),
            .I(N__22671));
    Span4Mux_h I__3019 (
            .O(N__22680),
            .I(N__22668));
    Span4Mux_v I__3018 (
            .O(N__22677),
            .I(N__22661));
    LocalMux I__3017 (
            .O(N__22674),
            .I(N__22661));
    Span4Mux_h I__3016 (
            .O(N__22671),
            .I(N__22661));
    Odrv4 I__3015 (
            .O(N__22668),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__3014 (
            .O(N__22661),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__3013 (
            .O(N__22656),
            .I(N__22653));
    LocalMux I__3012 (
            .O(N__22653),
            .I(N__22650));
    Odrv4 I__3011 (
            .O(N__22650),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ));
    CascadeMux I__3010 (
            .O(N__22647),
            .I(N__22644));
    InMux I__3009 (
            .O(N__22644),
            .I(N__22640));
    InMux I__3008 (
            .O(N__22643),
            .I(N__22637));
    LocalMux I__3007 (
            .O(N__22640),
            .I(N__22632));
    LocalMux I__3006 (
            .O(N__22637),
            .I(N__22632));
    Span4Mux_v I__3005 (
            .O(N__22632),
            .I(N__22627));
    InMux I__3004 (
            .O(N__22631),
            .I(N__22622));
    InMux I__3003 (
            .O(N__22630),
            .I(N__22622));
    Odrv4 I__3002 (
            .O(N__22627),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__3001 (
            .O(N__22622),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__3000 (
            .O(N__22617),
            .I(N__22614));
    LocalMux I__2999 (
            .O(N__22614),
            .I(N__22609));
    InMux I__2998 (
            .O(N__22613),
            .I(N__22606));
    CascadeMux I__2997 (
            .O(N__22612),
            .I(N__22603));
    Span4Mux_v I__2996 (
            .O(N__22609),
            .I(N__22597));
    LocalMux I__2995 (
            .O(N__22606),
            .I(N__22597));
    InMux I__2994 (
            .O(N__22603),
            .I(N__22592));
    InMux I__2993 (
            .O(N__22602),
            .I(N__22592));
    Odrv4 I__2992 (
            .O(N__22597),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__2991 (
            .O(N__22592),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__2990 (
            .O(N__22587),
            .I(\current_shift_inst.PI_CTRL.N_46_21_cascade_ ));
    InMux I__2989 (
            .O(N__22584),
            .I(N__22581));
    LocalMux I__2988 (
            .O(N__22581),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ));
    InMux I__2987 (
            .O(N__22578),
            .I(N__22575));
    LocalMux I__2986 (
            .O(N__22575),
            .I(N__22572));
    Span4Mux_v I__2985 (
            .O(N__22572),
            .I(N__22569));
    Odrv4 I__2984 (
            .O(N__22569),
            .I(\current_shift_inst.PI_CTRL.N_34 ));
    InMux I__2983 (
            .O(N__22566),
            .I(N__22561));
    InMux I__2982 (
            .O(N__22565),
            .I(N__22557));
    InMux I__2981 (
            .O(N__22564),
            .I(N__22554));
    LocalMux I__2980 (
            .O(N__22561),
            .I(N__22551));
    InMux I__2979 (
            .O(N__22560),
            .I(N__22548));
    LocalMux I__2978 (
            .O(N__22557),
            .I(N__22543));
    LocalMux I__2977 (
            .O(N__22554),
            .I(N__22543));
    Odrv12 I__2976 (
            .O(N__22551),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__2975 (
            .O(N__22548),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv12 I__2974 (
            .O(N__22543),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__2973 (
            .O(N__22536),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__2972 (
            .O(N__22533),
            .I(N__22530));
    LocalMux I__2971 (
            .O(N__22530),
            .I(N__22524));
    InMux I__2970 (
            .O(N__22529),
            .I(N__22521));
    CascadeMux I__2969 (
            .O(N__22528),
            .I(N__22518));
    InMux I__2968 (
            .O(N__22527),
            .I(N__22515));
    Span4Mux_v I__2967 (
            .O(N__22524),
            .I(N__22510));
    LocalMux I__2966 (
            .O(N__22521),
            .I(N__22510));
    InMux I__2965 (
            .O(N__22518),
            .I(N__22507));
    LocalMux I__2964 (
            .O(N__22515),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__2963 (
            .O(N__22510),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__2962 (
            .O(N__22507),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__2961 (
            .O(N__22500),
            .I(N__22497));
    LocalMux I__2960 (
            .O(N__22497),
            .I(\current_shift_inst.PI_CTRL.N_44 ));
    CascadeMux I__2959 (
            .O(N__22494),
            .I(\current_shift_inst.PI_CTRL.N_44_cascade_ ));
    InMux I__2958 (
            .O(N__22491),
            .I(N__22486));
    InMux I__2957 (
            .O(N__22490),
            .I(N__22480));
    InMux I__2956 (
            .O(N__22489),
            .I(N__22480));
    LocalMux I__2955 (
            .O(N__22486),
            .I(N__22477));
    InMux I__2954 (
            .O(N__22485),
            .I(N__22474));
    LocalMux I__2953 (
            .O(N__22480),
            .I(N__22471));
    Odrv12 I__2952 (
            .O(N__22477),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__2951 (
            .O(N__22474),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__2950 (
            .O(N__22471),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    CascadeMux I__2949 (
            .O(N__22464),
            .I(N__22461));
    InMux I__2948 (
            .O(N__22461),
            .I(N__22458));
    LocalMux I__2947 (
            .O(N__22458),
            .I(N__22452));
    InMux I__2946 (
            .O(N__22457),
            .I(N__22447));
    InMux I__2945 (
            .O(N__22456),
            .I(N__22447));
    InMux I__2944 (
            .O(N__22455),
            .I(N__22444));
    Span4Mux_v I__2943 (
            .O(N__22452),
            .I(N__22439));
    LocalMux I__2942 (
            .O(N__22447),
            .I(N__22439));
    LocalMux I__2941 (
            .O(N__22444),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__2940 (
            .O(N__22439),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    CascadeMux I__2939 (
            .O(N__22434),
            .I(N__22429));
    InMux I__2938 (
            .O(N__22433),
            .I(N__22426));
    InMux I__2937 (
            .O(N__22432),
            .I(N__22420));
    InMux I__2936 (
            .O(N__22429),
            .I(N__22420));
    LocalMux I__2935 (
            .O(N__22426),
            .I(N__22417));
    InMux I__2934 (
            .O(N__22425),
            .I(N__22414));
    LocalMux I__2933 (
            .O(N__22420),
            .I(N__22411));
    Odrv4 I__2932 (
            .O(N__22417),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__2931 (
            .O(N__22414),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__2930 (
            .O(N__22411),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__2929 (
            .O(N__22404),
            .I(N__22399));
    InMux I__2928 (
            .O(N__22403),
            .I(N__22393));
    InMux I__2927 (
            .O(N__22402),
            .I(N__22393));
    LocalMux I__2926 (
            .O(N__22399),
            .I(N__22390));
    InMux I__2925 (
            .O(N__22398),
            .I(N__22387));
    LocalMux I__2924 (
            .O(N__22393),
            .I(N__22384));
    Odrv4 I__2923 (
            .O(N__22390),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__2922 (
            .O(N__22387),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__2921 (
            .O(N__22384),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__2920 (
            .O(N__22377),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ));
    CascadeMux I__2919 (
            .O(N__22374),
            .I(N__22371));
    InMux I__2918 (
            .O(N__22371),
            .I(N__22368));
    LocalMux I__2917 (
            .O(N__22368),
            .I(N__22363));
    InMux I__2916 (
            .O(N__22367),
            .I(N__22358));
    InMux I__2915 (
            .O(N__22366),
            .I(N__22358));
    Span4Mux_v I__2914 (
            .O(N__22363),
            .I(N__22352));
    LocalMux I__2913 (
            .O(N__22358),
            .I(N__22352));
    InMux I__2912 (
            .O(N__22357),
            .I(N__22349));
    Odrv4 I__2911 (
            .O(N__22352),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__2910 (
            .O(N__22349),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__2909 (
            .O(N__22344),
            .I(N__22341));
    LocalMux I__2908 (
            .O(N__22341),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ));
    CascadeMux I__2907 (
            .O(N__22338),
            .I(clk_10khz_RNIIENAZ0Z2_cascade_));
    InMux I__2906 (
            .O(N__22335),
            .I(N__22332));
    LocalMux I__2905 (
            .O(N__22332),
            .I(clk_10khz_RNIIENAZ0Z2));
    InMux I__2904 (
            .O(N__22329),
            .I(N__22325));
    InMux I__2903 (
            .O(N__22328),
            .I(N__22322));
    LocalMux I__2902 (
            .O(N__22325),
            .I(N__22318));
    LocalMux I__2901 (
            .O(N__22322),
            .I(N__22315));
    InMux I__2900 (
            .O(N__22321),
            .I(N__22309));
    Span4Mux_v I__2899 (
            .O(N__22318),
            .I(N__22304));
    Span4Mux_v I__2898 (
            .O(N__22315),
            .I(N__22304));
    InMux I__2897 (
            .O(N__22314),
            .I(N__22301));
    InMux I__2896 (
            .O(N__22313),
            .I(N__22296));
    InMux I__2895 (
            .O(N__22312),
            .I(N__22296));
    LocalMux I__2894 (
            .O(N__22309),
            .I(N__22293));
    Odrv4 I__2893 (
            .O(N__22304),
            .I(un2_counter_8));
    LocalMux I__2892 (
            .O(N__22301),
            .I(un2_counter_8));
    LocalMux I__2891 (
            .O(N__22296),
            .I(un2_counter_8));
    Odrv4 I__2890 (
            .O(N__22293),
            .I(un2_counter_8));
    CascadeMux I__2889 (
            .O(N__22284),
            .I(N__22280));
    InMux I__2888 (
            .O(N__22283),
            .I(N__22277));
    InMux I__2887 (
            .O(N__22280),
            .I(N__22274));
    LocalMux I__2886 (
            .O(N__22277),
            .I(N__22267));
    LocalMux I__2885 (
            .O(N__22274),
            .I(N__22264));
    InMux I__2884 (
            .O(N__22273),
            .I(N__22261));
    InMux I__2883 (
            .O(N__22272),
            .I(N__22258));
    InMux I__2882 (
            .O(N__22271),
            .I(N__22253));
    InMux I__2881 (
            .O(N__22270),
            .I(N__22253));
    Span4Mux_v I__2880 (
            .O(N__22267),
            .I(N__22248));
    Span4Mux_v I__2879 (
            .O(N__22264),
            .I(N__22248));
    LocalMux I__2878 (
            .O(N__22261),
            .I(N__22245));
    LocalMux I__2877 (
            .O(N__22258),
            .I(un2_counter_7));
    LocalMux I__2876 (
            .O(N__22253),
            .I(un2_counter_7));
    Odrv4 I__2875 (
            .O(N__22248),
            .I(un2_counter_7));
    Odrv4 I__2874 (
            .O(N__22245),
            .I(un2_counter_7));
    InMux I__2873 (
            .O(N__22236),
            .I(N__22232));
    InMux I__2872 (
            .O(N__22235),
            .I(N__22229));
    LocalMux I__2871 (
            .O(N__22232),
            .I(N__22222));
    LocalMux I__2870 (
            .O(N__22229),
            .I(N__22219));
    InMux I__2869 (
            .O(N__22228),
            .I(N__22216));
    InMux I__2868 (
            .O(N__22227),
            .I(N__22213));
    InMux I__2867 (
            .O(N__22226),
            .I(N__22208));
    InMux I__2866 (
            .O(N__22225),
            .I(N__22208));
    Span4Mux_v I__2865 (
            .O(N__22222),
            .I(N__22201));
    Span4Mux_v I__2864 (
            .O(N__22219),
            .I(N__22201));
    LocalMux I__2863 (
            .O(N__22216),
            .I(N__22201));
    LocalMux I__2862 (
            .O(N__22213),
            .I(un2_counter_9));
    LocalMux I__2861 (
            .O(N__22208),
            .I(un2_counter_9));
    Odrv4 I__2860 (
            .O(N__22201),
            .I(un2_counter_9));
    CascadeMux I__2859 (
            .O(N__22194),
            .I(N__22188));
    InMux I__2858 (
            .O(N__22193),
            .I(N__22183));
    InMux I__2857 (
            .O(N__22192),
            .I(N__22183));
    InMux I__2856 (
            .O(N__22191),
            .I(N__22178));
    InMux I__2855 (
            .O(N__22188),
            .I(N__22178));
    LocalMux I__2854 (
            .O(N__22183),
            .I(clk_10khz_i));
    LocalMux I__2853 (
            .O(N__22178),
            .I(clk_10khz_i));
    InMux I__2852 (
            .O(N__22173),
            .I(N__22170));
    LocalMux I__2851 (
            .O(N__22170),
            .I(N__22167));
    Odrv4 I__2850 (
            .O(N__22167),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    CascadeMux I__2849 (
            .O(N__22164),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    CascadeMux I__2848 (
            .O(N__22161),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__2847 (
            .O(N__22158),
            .I(N__22155));
    LocalMux I__2846 (
            .O(N__22155),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    CascadeMux I__2845 (
            .O(N__22152),
            .I(N__22149));
    InMux I__2844 (
            .O(N__22149),
            .I(N__22146));
    LocalMux I__2843 (
            .O(N__22146),
            .I(N__22143));
    Span4Mux_h I__2842 (
            .O(N__22143),
            .I(N__22140));
    Odrv4 I__2841 (
            .O(N__22140),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__2840 (
            .O(N__22137),
            .I(N__22134));
    InMux I__2839 (
            .O(N__22134),
            .I(N__22131));
    LocalMux I__2838 (
            .O(N__22131),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    CascadeMux I__2837 (
            .O(N__22128),
            .I(N__22125));
    InMux I__2836 (
            .O(N__22125),
            .I(N__22122));
    LocalMux I__2835 (
            .O(N__22122),
            .I(N__22119));
    Span4Mux_h I__2834 (
            .O(N__22119),
            .I(N__22116));
    Odrv4 I__2833 (
            .O(N__22116),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__2832 (
            .O(N__22113),
            .I(N__22110));
    InMux I__2831 (
            .O(N__22110),
            .I(N__22107));
    LocalMux I__2830 (
            .O(N__22107),
            .I(N__22104));
    Odrv4 I__2829 (
            .O(N__22104),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__2828 (
            .O(N__22101),
            .I(N__22098));
    InMux I__2827 (
            .O(N__22098),
            .I(N__22095));
    LocalMux I__2826 (
            .O(N__22095),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    CascadeMux I__2825 (
            .O(N__22092),
            .I(N__22089));
    InMux I__2824 (
            .O(N__22089),
            .I(N__22086));
    LocalMux I__2823 (
            .O(N__22086),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    InMux I__2822 (
            .O(N__22083),
            .I(N__22080));
    LocalMux I__2821 (
            .O(N__22080),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    CascadeMux I__2820 (
            .O(N__22077),
            .I(N__22074));
    InMux I__2819 (
            .O(N__22074),
            .I(N__22068));
    InMux I__2818 (
            .O(N__22073),
            .I(N__22065));
    InMux I__2817 (
            .O(N__22072),
            .I(N__22062));
    CascadeMux I__2816 (
            .O(N__22071),
            .I(N__22059));
    LocalMux I__2815 (
            .O(N__22068),
            .I(N__22054));
    LocalMux I__2814 (
            .O(N__22065),
            .I(N__22054));
    LocalMux I__2813 (
            .O(N__22062),
            .I(N__22051));
    InMux I__2812 (
            .O(N__22059),
            .I(N__22048));
    Span4Mux_h I__2811 (
            .O(N__22054),
            .I(N__22045));
    Odrv4 I__2810 (
            .O(N__22051),
            .I(counterZ0Z_0));
    LocalMux I__2809 (
            .O(N__22048),
            .I(counterZ0Z_0));
    Odrv4 I__2808 (
            .O(N__22045),
            .I(counterZ0Z_0));
    InMux I__2807 (
            .O(N__22038),
            .I(N__22035));
    LocalMux I__2806 (
            .O(N__22035),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__2805 (
            .O(N__22032),
            .I(N__22029));
    InMux I__2804 (
            .O(N__22029),
            .I(N__22026));
    LocalMux I__2803 (
            .O(N__22026),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__2802 (
            .O(N__22023),
            .I(N__22020));
    InMux I__2801 (
            .O(N__22020),
            .I(N__22017));
    LocalMux I__2800 (
            .O(N__22017),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__2799 (
            .O(N__22014),
            .I(N__22011));
    LocalMux I__2798 (
            .O(N__22011),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    CascadeMux I__2797 (
            .O(N__22008),
            .I(N__22005));
    InMux I__2796 (
            .O(N__22005),
            .I(N__22002));
    LocalMux I__2795 (
            .O(N__22002),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    InMux I__2794 (
            .O(N__21999),
            .I(N__21996));
    LocalMux I__2793 (
            .O(N__21996),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    CascadeMux I__2792 (
            .O(N__21993),
            .I(N__21990));
    InMux I__2791 (
            .O(N__21990),
            .I(N__21987));
    LocalMux I__2790 (
            .O(N__21987),
            .I(N__21984));
    Odrv4 I__2789 (
            .O(N__21984),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    CascadeMux I__2788 (
            .O(N__21981),
            .I(N__21978));
    InMux I__2787 (
            .O(N__21978),
            .I(N__21975));
    LocalMux I__2786 (
            .O(N__21975),
            .I(N__21972));
    Odrv4 I__2785 (
            .O(N__21972),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    InMux I__2784 (
            .O(N__21969),
            .I(N__21966));
    LocalMux I__2783 (
            .O(N__21966),
            .I(N__21963));
    Odrv12 I__2782 (
            .O(N__21963),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    CascadeMux I__2781 (
            .O(N__21960),
            .I(N__21957));
    InMux I__2780 (
            .O(N__21957),
            .I(N__21954));
    LocalMux I__2779 (
            .O(N__21954),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    InMux I__2778 (
            .O(N__21951),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ));
    InMux I__2777 (
            .O(N__21948),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    InMux I__2776 (
            .O(N__21945),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    InMux I__2775 (
            .O(N__21942),
            .I(N__21939));
    LocalMux I__2774 (
            .O(N__21939),
            .I(N__21936));
    Odrv4 I__2773 (
            .O(N__21936),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__2772 (
            .O(N__21933),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    InMux I__2771 (
            .O(N__21930),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    InMux I__2770 (
            .O(N__21927),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__2769 (
            .O(N__21924),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    CascadeMux I__2768 (
            .O(N__21921),
            .I(N__21918));
    InMux I__2767 (
            .O(N__21918),
            .I(N__21915));
    LocalMux I__2766 (
            .O(N__21915),
            .I(N__21912));
    Odrv12 I__2765 (
            .O(N__21912),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__2764 (
            .O(N__21909),
            .I(N__21906));
    InMux I__2763 (
            .O(N__21906),
            .I(N__21903));
    LocalMux I__2762 (
            .O(N__21903),
            .I(N__21900));
    Odrv4 I__2761 (
            .O(N__21900),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__2760 (
            .O(N__21897),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ));
    InMux I__2759 (
            .O(N__21894),
            .I(N__21891));
    LocalMux I__2758 (
            .O(N__21891),
            .I(N__21888));
    Odrv4 I__2757 (
            .O(N__21888),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__2756 (
            .O(N__21885),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    InMux I__2755 (
            .O(N__21882),
            .I(N__21879));
    LocalMux I__2754 (
            .O(N__21879),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__2753 (
            .O(N__21876),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    CascadeMux I__2752 (
            .O(N__21873),
            .I(N__21870));
    InMux I__2751 (
            .O(N__21870),
            .I(N__21867));
    LocalMux I__2750 (
            .O(N__21867),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__2749 (
            .O(N__21864),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    InMux I__2748 (
            .O(N__21861),
            .I(N__21858));
    LocalMux I__2747 (
            .O(N__21858),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__2746 (
            .O(N__21855),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__2745 (
            .O(N__21852),
            .I(N__21849));
    InMux I__2744 (
            .O(N__21849),
            .I(N__21846));
    LocalMux I__2743 (
            .O(N__21846),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__2742 (
            .O(N__21843),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    InMux I__2741 (
            .O(N__21840),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    InMux I__2740 (
            .O(N__21837),
            .I(bfn_5_13_0_));
    InMux I__2739 (
            .O(N__21834),
            .I(N__21831));
    LocalMux I__2738 (
            .O(N__21831),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__2737 (
            .O(N__21828),
            .I(bfn_5_11_0_));
    CascadeMux I__2736 (
            .O(N__21825),
            .I(N__21822));
    InMux I__2735 (
            .O(N__21822),
            .I(N__21819));
    LocalMux I__2734 (
            .O(N__21819),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__2733 (
            .O(N__21816),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ));
    InMux I__2732 (
            .O(N__21813),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    InMux I__2731 (
            .O(N__21810),
            .I(N__21807));
    LocalMux I__2730 (
            .O(N__21807),
            .I(N__21804));
    Odrv4 I__2729 (
            .O(N__21804),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__2728 (
            .O(N__21801),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    InMux I__2727 (
            .O(N__21798),
            .I(N__21795));
    LocalMux I__2726 (
            .O(N__21795),
            .I(N__21792));
    Odrv4 I__2725 (
            .O(N__21792),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__2724 (
            .O(N__21789),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__2723 (
            .O(N__21786),
            .I(N__21783));
    InMux I__2722 (
            .O(N__21783),
            .I(N__21780));
    LocalMux I__2721 (
            .O(N__21780),
            .I(N__21777));
    Odrv4 I__2720 (
            .O(N__21777),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__2719 (
            .O(N__21774),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    InMux I__2718 (
            .O(N__21771),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    InMux I__2717 (
            .O(N__21768),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    InMux I__2716 (
            .O(N__21765),
            .I(N__21762));
    LocalMux I__2715 (
            .O(N__21762),
            .I(N__21759));
    Odrv4 I__2714 (
            .O(N__21759),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__2713 (
            .O(N__21756),
            .I(bfn_5_12_0_));
    InMux I__2712 (
            .O(N__21753),
            .I(N__21750));
    LocalMux I__2711 (
            .O(N__21750),
            .I(N__21747));
    Span4Mux_v I__2710 (
            .O(N__21747),
            .I(N__21742));
    InMux I__2709 (
            .O(N__21746),
            .I(N__21739));
    InMux I__2708 (
            .O(N__21745),
            .I(N__21736));
    Odrv4 I__2707 (
            .O(N__21742),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__2706 (
            .O(N__21739),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__2705 (
            .O(N__21736),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__2704 (
            .O(N__21729),
            .I(N__21726));
    LocalMux I__2703 (
            .O(N__21726),
            .I(N__21723));
    Span4Mux_v I__2702 (
            .O(N__21723),
            .I(N__21718));
    InMux I__2701 (
            .O(N__21722),
            .I(N__21715));
    InMux I__2700 (
            .O(N__21721),
            .I(N__21712));
    Odrv4 I__2699 (
            .O(N__21718),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__2698 (
            .O(N__21715),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__2697 (
            .O(N__21712),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__2696 (
            .O(N__21705),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ));
    CascadeMux I__2695 (
            .O(N__21702),
            .I(N__21699));
    InMux I__2694 (
            .O(N__21699),
            .I(N__21694));
    InMux I__2693 (
            .O(N__21698),
            .I(N__21691));
    InMux I__2692 (
            .O(N__21697),
            .I(N__21688));
    LocalMux I__2691 (
            .O(N__21694),
            .I(N__21683));
    LocalMux I__2690 (
            .O(N__21691),
            .I(N__21683));
    LocalMux I__2689 (
            .O(N__21688),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__2688 (
            .O(N__21683),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__2687 (
            .O(N__21678),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    InMux I__2686 (
            .O(N__21675),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    InMux I__2685 (
            .O(N__21672),
            .I(N__21669));
    LocalMux I__2684 (
            .O(N__21669),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__2683 (
            .O(N__21666),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    InMux I__2682 (
            .O(N__21663),
            .I(N__21660));
    LocalMux I__2681 (
            .O(N__21660),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__2680 (
            .O(N__21657),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    InMux I__2679 (
            .O(N__21654),
            .I(N__21651));
    LocalMux I__2678 (
            .O(N__21651),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__2677 (
            .O(N__21648),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    InMux I__2676 (
            .O(N__21645),
            .I(N__21642));
    LocalMux I__2675 (
            .O(N__21642),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__2674 (
            .O(N__21639),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    InMux I__2673 (
            .O(N__21636),
            .I(N__21633));
    LocalMux I__2672 (
            .O(N__21633),
            .I(N__21630));
    Odrv4 I__2671 (
            .O(N__21630),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    InMux I__2670 (
            .O(N__21627),
            .I(N__21624));
    LocalMux I__2669 (
            .O(N__21624),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    InMux I__2668 (
            .O(N__21621),
            .I(N__21618));
    LocalMux I__2667 (
            .O(N__21618),
            .I(N__21615));
    Odrv4 I__2666 (
            .O(N__21615),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__2665 (
            .O(N__21612),
            .I(N__21609));
    LocalMux I__2664 (
            .O(N__21609),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    InMux I__2663 (
            .O(N__21606),
            .I(N__21603));
    LocalMux I__2662 (
            .O(N__21603),
            .I(N__21600));
    Span4Mux_v I__2661 (
            .O(N__21600),
            .I(N__21597));
    Odrv4 I__2660 (
            .O(N__21597),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__2659 (
            .O(N__21594),
            .I(N__21590));
    InMux I__2658 (
            .O(N__21593),
            .I(N__21587));
    LocalMux I__2657 (
            .O(N__21590),
            .I(counterZ0Z_2));
    LocalMux I__2656 (
            .O(N__21587),
            .I(counterZ0Z_2));
    InMux I__2655 (
            .O(N__21582),
            .I(N__21577));
    InMux I__2654 (
            .O(N__21581),
            .I(N__21574));
    InMux I__2653 (
            .O(N__21580),
            .I(N__21571));
    LocalMux I__2652 (
            .O(N__21577),
            .I(counterZ0Z_1));
    LocalMux I__2651 (
            .O(N__21574),
            .I(counterZ0Z_1));
    LocalMux I__2650 (
            .O(N__21571),
            .I(counterZ0Z_1));
    CascadeMux I__2649 (
            .O(N__21564),
            .I(un2_counter_5_cascade_));
    InMux I__2648 (
            .O(N__21561),
            .I(N__21557));
    InMux I__2647 (
            .O(N__21560),
            .I(N__21554));
    LocalMux I__2646 (
            .O(N__21557),
            .I(counterZ0Z_8));
    LocalMux I__2645 (
            .O(N__21554),
            .I(counterZ0Z_8));
    InMux I__2644 (
            .O(N__21549),
            .I(N__21545));
    InMux I__2643 (
            .O(N__21548),
            .I(N__21542));
    LocalMux I__2642 (
            .O(N__21545),
            .I(counterZ0Z_11));
    LocalMux I__2641 (
            .O(N__21542),
            .I(counterZ0Z_11));
    InMux I__2640 (
            .O(N__21537),
            .I(N__21533));
    InMux I__2639 (
            .O(N__21536),
            .I(N__21530));
    LocalMux I__2638 (
            .O(N__21533),
            .I(counterZ0Z_9));
    LocalMux I__2637 (
            .O(N__21530),
            .I(counterZ0Z_9));
    InMux I__2636 (
            .O(N__21525),
            .I(N__21521));
    InMux I__2635 (
            .O(N__21524),
            .I(N__21518));
    LocalMux I__2634 (
            .O(N__21521),
            .I(counterZ0Z_5));
    LocalMux I__2633 (
            .O(N__21518),
            .I(counterZ0Z_5));
    InMux I__2632 (
            .O(N__21513),
            .I(N__21509));
    InMux I__2631 (
            .O(N__21512),
            .I(N__21506));
    LocalMux I__2630 (
            .O(N__21509),
            .I(counterZ0Z_4));
    LocalMux I__2629 (
            .O(N__21506),
            .I(counterZ0Z_4));
    CascadeMux I__2628 (
            .O(N__21501),
            .I(N__21497));
    InMux I__2627 (
            .O(N__21500),
            .I(N__21494));
    InMux I__2626 (
            .O(N__21497),
            .I(N__21491));
    LocalMux I__2625 (
            .O(N__21494),
            .I(counterZ0Z_6));
    LocalMux I__2624 (
            .O(N__21491),
            .I(counterZ0Z_6));
    InMux I__2623 (
            .O(N__21486),
            .I(N__21482));
    InMux I__2622 (
            .O(N__21485),
            .I(N__21479));
    LocalMux I__2621 (
            .O(N__21482),
            .I(counterZ0Z_3));
    LocalMux I__2620 (
            .O(N__21479),
            .I(counterZ0Z_3));
    InMux I__2619 (
            .O(N__21474),
            .I(N__21471));
    LocalMux I__2618 (
            .O(N__21471),
            .I(N__21468));
    Span4Mux_h I__2617 (
            .O(N__21468),
            .I(N__21465));
    Odrv4 I__2616 (
            .O(N__21465),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__2615 (
            .O(N__21462),
            .I(N__21459));
    LocalMux I__2614 (
            .O(N__21459),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    InMux I__2613 (
            .O(N__21456),
            .I(N__21453));
    LocalMux I__2612 (
            .O(N__21453),
            .I(N__21450));
    Span4Mux_v I__2611 (
            .O(N__21450),
            .I(N__21447));
    Odrv4 I__2610 (
            .O(N__21447),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    CascadeMux I__2609 (
            .O(N__21444),
            .I(N__21441));
    InMux I__2608 (
            .O(N__21441),
            .I(N__21438));
    LocalMux I__2607 (
            .O(N__21438),
            .I(counter_RNO_0Z0Z_12));
    CascadeMux I__2606 (
            .O(N__21435),
            .I(N__21431));
    InMux I__2605 (
            .O(N__21434),
            .I(N__21428));
    InMux I__2604 (
            .O(N__21431),
            .I(N__21425));
    LocalMux I__2603 (
            .O(N__21428),
            .I(counterZ0Z_12));
    LocalMux I__2602 (
            .O(N__21425),
            .I(counterZ0Z_12));
    CascadeMux I__2601 (
            .O(N__21420),
            .I(N__21417));
    InMux I__2600 (
            .O(N__21417),
            .I(N__21414));
    LocalMux I__2599 (
            .O(N__21414),
            .I(counter_RNO_0Z0Z_10));
    InMux I__2598 (
            .O(N__21411),
            .I(N__21407));
    InMux I__2597 (
            .O(N__21410),
            .I(N__21404));
    LocalMux I__2596 (
            .O(N__21407),
            .I(counterZ0Z_10));
    LocalMux I__2595 (
            .O(N__21404),
            .I(counterZ0Z_10));
    InMux I__2594 (
            .O(N__21399),
            .I(N__21393));
    InMux I__2593 (
            .O(N__21398),
            .I(N__21393));
    LocalMux I__2592 (
            .O(N__21393),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2591 (
            .O(N__21390),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2590 (
            .O(N__21387),
            .I(N__21383));
    InMux I__2589 (
            .O(N__21386),
            .I(N__21380));
    LocalMux I__2588 (
            .O(N__21383),
            .I(N__21375));
    LocalMux I__2587 (
            .O(N__21380),
            .I(N__21375));
    Span4Mux_v I__2586 (
            .O(N__21375),
            .I(N__21372));
    Odrv4 I__2585 (
            .O(N__21372),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2584 (
            .O(N__21369),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2583 (
            .O(N__21366),
            .I(N__21360));
    InMux I__2582 (
            .O(N__21365),
            .I(N__21360));
    LocalMux I__2581 (
            .O(N__21360),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2580 (
            .O(N__21357),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2579 (
            .O(N__21354),
            .I(N__21351));
    LocalMux I__2578 (
            .O(N__21351),
            .I(N__21347));
    CascadeMux I__2577 (
            .O(N__21350),
            .I(N__21344));
    Span4Mux_h I__2576 (
            .O(N__21347),
            .I(N__21341));
    InMux I__2575 (
            .O(N__21344),
            .I(N__21338));
    Odrv4 I__2574 (
            .O(N__21341),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__2573 (
            .O(N__21338),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2572 (
            .O(N__21333),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    CascadeMux I__2571 (
            .O(N__21330),
            .I(N__21327));
    InMux I__2570 (
            .O(N__21327),
            .I(N__21324));
    LocalMux I__2569 (
            .O(N__21324),
            .I(N__21320));
    InMux I__2568 (
            .O(N__21323),
            .I(N__21317));
    Span4Mux_h I__2567 (
            .O(N__21320),
            .I(N__21314));
    LocalMux I__2566 (
            .O(N__21317),
            .I(N__21311));
    Odrv4 I__2565 (
            .O(N__21314),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    Odrv4 I__2564 (
            .O(N__21311),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2563 (
            .O(N__21306),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2562 (
            .O(N__21303),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2561 (
            .O(N__21300),
            .I(N__21297));
    LocalMux I__2560 (
            .O(N__21297),
            .I(N__21288));
    InMux I__2559 (
            .O(N__21296),
            .I(N__21285));
    InMux I__2558 (
            .O(N__21295),
            .I(N__21281));
    InMux I__2557 (
            .O(N__21294),
            .I(N__21272));
    InMux I__2556 (
            .O(N__21293),
            .I(N__21272));
    InMux I__2555 (
            .O(N__21292),
            .I(N__21272));
    InMux I__2554 (
            .O(N__21291),
            .I(N__21272));
    Span4Mux_v I__2553 (
            .O(N__21288),
            .I(N__21267));
    LocalMux I__2552 (
            .O(N__21285),
            .I(N__21267));
    CascadeMux I__2551 (
            .O(N__21284),
            .I(N__21262));
    LocalMux I__2550 (
            .O(N__21281),
            .I(N__21259));
    LocalMux I__2549 (
            .O(N__21272),
            .I(N__21254));
    Span4Mux_h I__2548 (
            .O(N__21267),
            .I(N__21254));
    InMux I__2547 (
            .O(N__21266),
            .I(N__21251));
    InMux I__2546 (
            .O(N__21265),
            .I(N__21246));
    InMux I__2545 (
            .O(N__21262),
            .I(N__21246));
    Span4Mux_v I__2544 (
            .O(N__21259),
            .I(N__21239));
    Span4Mux_v I__2543 (
            .O(N__21254),
            .I(N__21239));
    LocalMux I__2542 (
            .O(N__21251),
            .I(N__21239));
    LocalMux I__2541 (
            .O(N__21246),
            .I(N__21234));
    Span4Mux_h I__2540 (
            .O(N__21239),
            .I(N__21234));
    Span4Mux_v I__2539 (
            .O(N__21234),
            .I(N__21231));
    Odrv4 I__2538 (
            .O(N__21231),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__2537 (
            .O(N__21228),
            .I(N__21225));
    InMux I__2536 (
            .O(N__21225),
            .I(N__21222));
    LocalMux I__2535 (
            .O(N__21222),
            .I(counter_RNO_0Z0Z_7));
    InMux I__2534 (
            .O(N__21219),
            .I(N__21215));
    InMux I__2533 (
            .O(N__21218),
            .I(N__21212));
    LocalMux I__2532 (
            .O(N__21215),
            .I(counterZ0Z_7));
    LocalMux I__2531 (
            .O(N__21212),
            .I(counterZ0Z_7));
    InMux I__2530 (
            .O(N__21207),
            .I(N__21201));
    InMux I__2529 (
            .O(N__21206),
            .I(N__21201));
    LocalMux I__2528 (
            .O(N__21201),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2527 (
            .O(N__21198),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    InMux I__2526 (
            .O(N__21195),
            .I(N__21189));
    InMux I__2525 (
            .O(N__21194),
            .I(N__21189));
    LocalMux I__2524 (
            .O(N__21189),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2523 (
            .O(N__21186),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2522 (
            .O(N__21183),
            .I(N__21177));
    InMux I__2521 (
            .O(N__21182),
            .I(N__21177));
    LocalMux I__2520 (
            .O(N__21177),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2519 (
            .O(N__21174),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2518 (
            .O(N__21171),
            .I(N__21165));
    InMux I__2517 (
            .O(N__21170),
            .I(N__21165));
    LocalMux I__2516 (
            .O(N__21165),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2515 (
            .O(N__21162),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__2514 (
            .O(N__21159),
            .I(N__21156));
    InMux I__2513 (
            .O(N__21156),
            .I(N__21150));
    InMux I__2512 (
            .O(N__21155),
            .I(N__21150));
    LocalMux I__2511 (
            .O(N__21150),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2510 (
            .O(N__21147),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2509 (
            .O(N__21144),
            .I(N__21141));
    LocalMux I__2508 (
            .O(N__21141),
            .I(N__21137));
    InMux I__2507 (
            .O(N__21140),
            .I(N__21134));
    Odrv4 I__2506 (
            .O(N__21137),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    LocalMux I__2505 (
            .O(N__21134),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2504 (
            .O(N__21129),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2503 (
            .O(N__21126),
            .I(N__21122));
    CascadeMux I__2502 (
            .O(N__21125),
            .I(N__21119));
    LocalMux I__2501 (
            .O(N__21122),
            .I(N__21116));
    InMux I__2500 (
            .O(N__21119),
            .I(N__21113));
    Odrv4 I__2499 (
            .O(N__21116),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    LocalMux I__2498 (
            .O(N__21113),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2497 (
            .O(N__21108),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    CascadeMux I__2496 (
            .O(N__21105),
            .I(N__21102));
    InMux I__2495 (
            .O(N__21102),
            .I(N__21098));
    InMux I__2494 (
            .O(N__21101),
            .I(N__21095));
    LocalMux I__2493 (
            .O(N__21098),
            .I(N__21090));
    LocalMux I__2492 (
            .O(N__21095),
            .I(N__21090));
    Span4Mux_v I__2491 (
            .O(N__21090),
            .I(N__21087));
    Odrv4 I__2490 (
            .O(N__21087),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2489 (
            .O(N__21084),
            .I(bfn_4_16_0_));
    InMux I__2488 (
            .O(N__21081),
            .I(N__21077));
    InMux I__2487 (
            .O(N__21080),
            .I(N__21074));
    LocalMux I__2486 (
            .O(N__21077),
            .I(N__21071));
    LocalMux I__2485 (
            .O(N__21074),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    Odrv4 I__2484 (
            .O(N__21071),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2483 (
            .O(N__21066),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    CascadeMux I__2482 (
            .O(N__21063),
            .I(N__21060));
    InMux I__2481 (
            .O(N__21060),
            .I(N__21056));
    InMux I__2480 (
            .O(N__21059),
            .I(N__21052));
    LocalMux I__2479 (
            .O(N__21056),
            .I(N__21049));
    InMux I__2478 (
            .O(N__21055),
            .I(N__21046));
    LocalMux I__2477 (
            .O(N__21052),
            .I(N__21043));
    Span4Mux_v I__2476 (
            .O(N__21049),
            .I(N__21036));
    LocalMux I__2475 (
            .O(N__21046),
            .I(N__21036));
    Span4Mux_v I__2474 (
            .O(N__21043),
            .I(N__21036));
    Odrv4 I__2473 (
            .O(N__21036),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2472 (
            .O(N__21033),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    InMux I__2471 (
            .O(N__21030),
            .I(N__21027));
    LocalMux I__2470 (
            .O(N__21027),
            .I(N__21024));
    Span4Mux_h I__2469 (
            .O(N__21024),
            .I(N__21020));
    InMux I__2468 (
            .O(N__21023),
            .I(N__21017));
    Odrv4 I__2467 (
            .O(N__21020),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    LocalMux I__2466 (
            .O(N__21017),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2465 (
            .O(N__21012),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    CascadeMux I__2464 (
            .O(N__21009),
            .I(N__21006));
    InMux I__2463 (
            .O(N__21006),
            .I(N__21000));
    InMux I__2462 (
            .O(N__21005),
            .I(N__21000));
    LocalMux I__2461 (
            .O(N__21000),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2460 (
            .O(N__20997),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2459 (
            .O(N__20994),
            .I(N__20988));
    InMux I__2458 (
            .O(N__20993),
            .I(N__20988));
    LocalMux I__2457 (
            .O(N__20988),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2456 (
            .O(N__20985),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    CascadeMux I__2455 (
            .O(N__20982),
            .I(N__20978));
    InMux I__2454 (
            .O(N__20981),
            .I(N__20975));
    InMux I__2453 (
            .O(N__20978),
            .I(N__20972));
    LocalMux I__2452 (
            .O(N__20975),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    LocalMux I__2451 (
            .O(N__20972),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2450 (
            .O(N__20967),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2449 (
            .O(N__20964),
            .I(N__20961));
    LocalMux I__2448 (
            .O(N__20961),
            .I(N__20957));
    InMux I__2447 (
            .O(N__20960),
            .I(N__20954));
    Odrv4 I__2446 (
            .O(N__20957),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    LocalMux I__2445 (
            .O(N__20954),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2444 (
            .O(N__20949),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2443 (
            .O(N__20946),
            .I(N__20943));
    LocalMux I__2442 (
            .O(N__20943),
            .I(N__20940));
    Span4Mux_h I__2441 (
            .O(N__20940),
            .I(N__20936));
    InMux I__2440 (
            .O(N__20939),
            .I(N__20933));
    Odrv4 I__2439 (
            .O(N__20936),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2438 (
            .O(N__20933),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2437 (
            .O(N__20928),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__2436 (
            .O(N__20925),
            .I(N__20921));
    InMux I__2435 (
            .O(N__20924),
            .I(N__20918));
    LocalMux I__2434 (
            .O(N__20921),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    LocalMux I__2433 (
            .O(N__20918),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2432 (
            .O(N__20913),
            .I(bfn_4_15_0_));
    CascadeMux I__2431 (
            .O(N__20910),
            .I(N__20907));
    InMux I__2430 (
            .O(N__20907),
            .I(N__20904));
    LocalMux I__2429 (
            .O(N__20904),
            .I(N__20901));
    Odrv12 I__2428 (
            .O(N__20901),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__2427 (
            .O(N__20898),
            .I(N__20895));
    InMux I__2426 (
            .O(N__20895),
            .I(N__20892));
    LocalMux I__2425 (
            .O(N__20892),
            .I(N__20889));
    Span4Mux_v I__2424 (
            .O(N__20889),
            .I(N__20886));
    Span4Mux_h I__2423 (
            .O(N__20886),
            .I(N__20883));
    Odrv4 I__2422 (
            .O(N__20883),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2421 (
            .O(N__20880),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    InMux I__2420 (
            .O(N__20877),
            .I(N__20874));
    LocalMux I__2419 (
            .O(N__20874),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__2418 (
            .O(N__20871),
            .I(N__20868));
    InMux I__2417 (
            .O(N__20868),
            .I(N__20865));
    LocalMux I__2416 (
            .O(N__20865),
            .I(N__20862));
    Span4Mux_h I__2415 (
            .O(N__20862),
            .I(N__20859));
    Span4Mux_v I__2414 (
            .O(N__20859),
            .I(N__20856));
    Odrv4 I__2413 (
            .O(N__20856),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2412 (
            .O(N__20853),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    CascadeMux I__2411 (
            .O(N__20850),
            .I(N__20847));
    InMux I__2410 (
            .O(N__20847),
            .I(N__20843));
    CascadeMux I__2409 (
            .O(N__20846),
            .I(N__20840));
    LocalMux I__2408 (
            .O(N__20843),
            .I(N__20837));
    InMux I__2407 (
            .O(N__20840),
            .I(N__20833));
    Span4Mux_h I__2406 (
            .O(N__20837),
            .I(N__20830));
    InMux I__2405 (
            .O(N__20836),
            .I(N__20827));
    LocalMux I__2404 (
            .O(N__20833),
            .I(N__20820));
    Span4Mux_v I__2403 (
            .O(N__20830),
            .I(N__20820));
    LocalMux I__2402 (
            .O(N__20827),
            .I(N__20820));
    Span4Mux_h I__2401 (
            .O(N__20820),
            .I(N__20817));
    Odrv4 I__2400 (
            .O(N__20817),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2399 (
            .O(N__20814),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    CascadeMux I__2398 (
            .O(N__20811),
            .I(N__20806));
    InMux I__2397 (
            .O(N__20810),
            .I(N__20800));
    InMux I__2396 (
            .O(N__20809),
            .I(N__20800));
    InMux I__2395 (
            .O(N__20806),
            .I(N__20797));
    InMux I__2394 (
            .O(N__20805),
            .I(N__20794));
    LocalMux I__2393 (
            .O(N__20800),
            .I(N__20791));
    LocalMux I__2392 (
            .O(N__20797),
            .I(N__20788));
    LocalMux I__2391 (
            .O(N__20794),
            .I(N__20785));
    Span4Mux_h I__2390 (
            .O(N__20791),
            .I(N__20782));
    Odrv4 I__2389 (
            .O(N__20788),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2388 (
            .O(N__20785),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2387 (
            .O(N__20782),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2386 (
            .O(N__20775),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2385 (
            .O(N__20772),
            .I(N__20769));
    LocalMux I__2384 (
            .O(N__20769),
            .I(N__20766));
    Odrv12 I__2383 (
            .O(N__20766),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__2382 (
            .O(N__20763),
            .I(N__20760));
    InMux I__2381 (
            .O(N__20760),
            .I(N__20757));
    LocalMux I__2380 (
            .O(N__20757),
            .I(N__20753));
    InMux I__2379 (
            .O(N__20756),
            .I(N__20750));
    Span4Mux_v I__2378 (
            .O(N__20753),
            .I(N__20744));
    LocalMux I__2377 (
            .O(N__20750),
            .I(N__20744));
    InMux I__2376 (
            .O(N__20749),
            .I(N__20741));
    Span4Mux_v I__2375 (
            .O(N__20744),
            .I(N__20736));
    LocalMux I__2374 (
            .O(N__20741),
            .I(N__20736));
    Odrv4 I__2373 (
            .O(N__20736),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2372 (
            .O(N__20733),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    CascadeMux I__2371 (
            .O(N__20730),
            .I(N__20727));
    InMux I__2370 (
            .O(N__20727),
            .I(N__20724));
    LocalMux I__2369 (
            .O(N__20724),
            .I(N__20719));
    InMux I__2368 (
            .O(N__20723),
            .I(N__20716));
    InMux I__2367 (
            .O(N__20722),
            .I(N__20713));
    Span4Mux_v I__2366 (
            .O(N__20719),
            .I(N__20708));
    LocalMux I__2365 (
            .O(N__20716),
            .I(N__20708));
    LocalMux I__2364 (
            .O(N__20713),
            .I(N__20705));
    Span4Mux_h I__2363 (
            .O(N__20708),
            .I(N__20702));
    Odrv4 I__2362 (
            .O(N__20705),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2361 (
            .O(N__20702),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2360 (
            .O(N__20697),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    CascadeMux I__2359 (
            .O(N__20694),
            .I(N__20691));
    InMux I__2358 (
            .O(N__20691),
            .I(N__20688));
    LocalMux I__2357 (
            .O(N__20688),
            .I(N__20685));
    Span4Mux_v I__2356 (
            .O(N__20685),
            .I(N__20682));
    Odrv4 I__2355 (
            .O(N__20682),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__2354 (
            .O(N__20679),
            .I(N__20676));
    InMux I__2353 (
            .O(N__20676),
            .I(N__20671));
    InMux I__2352 (
            .O(N__20675),
            .I(N__20668));
    InMux I__2351 (
            .O(N__20674),
            .I(N__20665));
    LocalMux I__2350 (
            .O(N__20671),
            .I(N__20662));
    LocalMux I__2349 (
            .O(N__20668),
            .I(N__20659));
    LocalMux I__2348 (
            .O(N__20665),
            .I(N__20656));
    Span4Mux_v I__2347 (
            .O(N__20662),
            .I(N__20653));
    Span4Mux_v I__2346 (
            .O(N__20659),
            .I(N__20648));
    Span4Mux_s3_h I__2345 (
            .O(N__20656),
            .I(N__20648));
    Odrv4 I__2344 (
            .O(N__20653),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2343 (
            .O(N__20648),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2342 (
            .O(N__20643),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    CascadeMux I__2341 (
            .O(N__20640),
            .I(N__20637));
    InMux I__2340 (
            .O(N__20637),
            .I(N__20634));
    LocalMux I__2339 (
            .O(N__20634),
            .I(N__20630));
    InMux I__2338 (
            .O(N__20633),
            .I(N__20627));
    Span4Mux_v I__2337 (
            .O(N__20630),
            .I(N__20623));
    LocalMux I__2336 (
            .O(N__20627),
            .I(N__20620));
    InMux I__2335 (
            .O(N__20626),
            .I(N__20617));
    Span4Mux_s2_h I__2334 (
            .O(N__20623),
            .I(N__20610));
    Span4Mux_v I__2333 (
            .O(N__20620),
            .I(N__20610));
    LocalMux I__2332 (
            .O(N__20617),
            .I(N__20610));
    Odrv4 I__2331 (
            .O(N__20610),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2330 (
            .O(N__20607),
            .I(bfn_4_14_0_));
    CascadeMux I__2329 (
            .O(N__20604),
            .I(N__20601));
    InMux I__2328 (
            .O(N__20601),
            .I(N__20598));
    LocalMux I__2327 (
            .O(N__20598),
            .I(N__20595));
    Odrv4 I__2326 (
            .O(N__20595),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    CascadeMux I__2325 (
            .O(N__20592),
            .I(N__20589));
    InMux I__2324 (
            .O(N__20589),
            .I(N__20586));
    LocalMux I__2323 (
            .O(N__20586),
            .I(N__20583));
    Span4Mux_v I__2322 (
            .O(N__20583),
            .I(N__20580));
    Span4Mux_h I__2321 (
            .O(N__20580),
            .I(N__20577));
    Odrv4 I__2320 (
            .O(N__20577),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    CascadeMux I__2319 (
            .O(N__20574),
            .I(N__20571));
    InMux I__2318 (
            .O(N__20571),
            .I(N__20568));
    LocalMux I__2317 (
            .O(N__20568),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__2316 (
            .O(N__20565),
            .I(N__20558));
    InMux I__2315 (
            .O(N__20564),
            .I(N__20558));
    CascadeMux I__2314 (
            .O(N__20563),
            .I(N__20555));
    LocalMux I__2313 (
            .O(N__20558),
            .I(N__20545));
    InMux I__2312 (
            .O(N__20555),
            .I(N__20542));
    InMux I__2311 (
            .O(N__20554),
            .I(N__20535));
    InMux I__2310 (
            .O(N__20553),
            .I(N__20535));
    InMux I__2309 (
            .O(N__20552),
            .I(N__20535));
    InMux I__2308 (
            .O(N__20551),
            .I(N__20526));
    InMux I__2307 (
            .O(N__20550),
            .I(N__20526));
    InMux I__2306 (
            .O(N__20549),
            .I(N__20526));
    InMux I__2305 (
            .O(N__20548),
            .I(N__20526));
    Span4Mux_v I__2304 (
            .O(N__20545),
            .I(N__20517));
    LocalMux I__2303 (
            .O(N__20542),
            .I(N__20517));
    LocalMux I__2302 (
            .O(N__20535),
            .I(N__20517));
    LocalMux I__2301 (
            .O(N__20526),
            .I(N__20517));
    Span4Mux_h I__2300 (
            .O(N__20517),
            .I(N__20514));
    Span4Mux_v I__2299 (
            .O(N__20514),
            .I(N__20510));
    InMux I__2298 (
            .O(N__20513),
            .I(N__20507));
    Odrv4 I__2297 (
            .O(N__20510),
            .I(pwm_duty_input_6));
    LocalMux I__2296 (
            .O(N__20507),
            .I(pwm_duty_input_6));
    InMux I__2295 (
            .O(N__20502),
            .I(N__20493));
    InMux I__2294 (
            .O(N__20501),
            .I(N__20493));
    CascadeMux I__2293 (
            .O(N__20500),
            .I(N__20486));
    CascadeMux I__2292 (
            .O(N__20499),
            .I(N__20483));
    CascadeMux I__2291 (
            .O(N__20498),
            .I(N__20479));
    LocalMux I__2290 (
            .O(N__20493),
            .I(N__20476));
    InMux I__2289 (
            .O(N__20492),
            .I(N__20467));
    InMux I__2288 (
            .O(N__20491),
            .I(N__20467));
    InMux I__2287 (
            .O(N__20490),
            .I(N__20467));
    InMux I__2286 (
            .O(N__20489),
            .I(N__20467));
    InMux I__2285 (
            .O(N__20486),
            .I(N__20458));
    InMux I__2284 (
            .O(N__20483),
            .I(N__20458));
    InMux I__2283 (
            .O(N__20482),
            .I(N__20458));
    InMux I__2282 (
            .O(N__20479),
            .I(N__20458));
    Span4Mux_v I__2281 (
            .O(N__20476),
            .I(N__20451));
    LocalMux I__2280 (
            .O(N__20467),
            .I(N__20451));
    LocalMux I__2279 (
            .O(N__20458),
            .I(N__20451));
    Odrv4 I__2278 (
            .O(N__20451),
            .I(i8_mux));
    CascadeMux I__2277 (
            .O(N__20448),
            .I(N__20441));
    CascadeMux I__2276 (
            .O(N__20447),
            .I(N__20437));
    CascadeMux I__2275 (
            .O(N__20446),
            .I(N__20431));
    CascadeMux I__2274 (
            .O(N__20445),
            .I(N__20428));
    CascadeMux I__2273 (
            .O(N__20444),
            .I(N__20425));
    InMux I__2272 (
            .O(N__20441),
            .I(N__20419));
    InMux I__2271 (
            .O(N__20440),
            .I(N__20419));
    InMux I__2270 (
            .O(N__20437),
            .I(N__20416));
    InMux I__2269 (
            .O(N__20436),
            .I(N__20409));
    InMux I__2268 (
            .O(N__20435),
            .I(N__20409));
    InMux I__2267 (
            .O(N__20434),
            .I(N__20409));
    InMux I__2266 (
            .O(N__20431),
            .I(N__20400));
    InMux I__2265 (
            .O(N__20428),
            .I(N__20400));
    InMux I__2264 (
            .O(N__20425),
            .I(N__20400));
    InMux I__2263 (
            .O(N__20424),
            .I(N__20400));
    LocalMux I__2262 (
            .O(N__20419),
            .I(N__20397));
    LocalMux I__2261 (
            .O(N__20416),
            .I(N__20390));
    LocalMux I__2260 (
            .O(N__20409),
            .I(N__20390));
    LocalMux I__2259 (
            .O(N__20400),
            .I(N__20390));
    Span4Mux_h I__2258 (
            .O(N__20397),
            .I(N__20387));
    Odrv4 I__2257 (
            .O(N__20390),
            .I(N_28_mux));
    Odrv4 I__2256 (
            .O(N__20387),
            .I(N_28_mux));
    InMux I__2255 (
            .O(N__20382),
            .I(N__20379));
    LocalMux I__2254 (
            .O(N__20379),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__2253 (
            .O(N__20376),
            .I(N__20373));
    LocalMux I__2252 (
            .O(N__20373),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    InMux I__2251 (
            .O(N__20370),
            .I(bfn_4_6_0_));
    InMux I__2250 (
            .O(N__20367),
            .I(un5_counter_cry_9));
    InMux I__2249 (
            .O(N__20364),
            .I(un5_counter_cry_10));
    InMux I__2248 (
            .O(N__20361),
            .I(un5_counter_cry_11));
    InMux I__2247 (
            .O(N__20358),
            .I(N__20355));
    LocalMux I__2246 (
            .O(N__20355),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    InMux I__2245 (
            .O(N__20352),
            .I(N__20349));
    LocalMux I__2244 (
            .O(N__20349),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__2243 (
            .O(N__20346),
            .I(N__20343));
    LocalMux I__2242 (
            .O(N__20343),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__2241 (
            .O(N__20340),
            .I(N__20337));
    LocalMux I__2240 (
            .O(N__20337),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__2239 (
            .O(N__20334),
            .I(N__20331));
    LocalMux I__2238 (
            .O(N__20331),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__2237 (
            .O(N__20328),
            .I(un5_counter_cry_1));
    InMux I__2236 (
            .O(N__20325),
            .I(un5_counter_cry_2));
    InMux I__2235 (
            .O(N__20322),
            .I(un5_counter_cry_3));
    InMux I__2234 (
            .O(N__20319),
            .I(un5_counter_cry_4));
    InMux I__2233 (
            .O(N__20316),
            .I(un5_counter_cry_5));
    InMux I__2232 (
            .O(N__20313),
            .I(un5_counter_cry_6));
    InMux I__2231 (
            .O(N__20310),
            .I(un5_counter_cry_7));
    CascadeMux I__2230 (
            .O(N__20307),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    CascadeMux I__2229 (
            .O(N__20304),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ));
    InMux I__2228 (
            .O(N__20301),
            .I(N__20287));
    InMux I__2227 (
            .O(N__20300),
            .I(N__20287));
    InMux I__2226 (
            .O(N__20299),
            .I(N__20287));
    InMux I__2225 (
            .O(N__20298),
            .I(N__20287));
    InMux I__2224 (
            .O(N__20297),
            .I(N__20282));
    InMux I__2223 (
            .O(N__20296),
            .I(N__20282));
    LocalMux I__2222 (
            .O(N__20287),
            .I(N__20279));
    LocalMux I__2221 (
            .O(N__20282),
            .I(N__20276));
    Span4Mux_s3_h I__2220 (
            .O(N__20279),
            .I(N__20272));
    Span4Mux_s3_h I__2219 (
            .O(N__20276),
            .I(N__20269));
    InMux I__2218 (
            .O(N__20275),
            .I(N__20266));
    Odrv4 I__2217 (
            .O(N__20272),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2216 (
            .O(N__20269),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    LocalMux I__2215 (
            .O(N__20266),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2214 (
            .O(N__20259),
            .I(N__20256));
    LocalMux I__2213 (
            .O(N__20256),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__2212 (
            .O(N__20253),
            .I(N__20250));
    LocalMux I__2211 (
            .O(N__20250),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__2210 (
            .O(N__20247),
            .I(N__20244));
    LocalMux I__2209 (
            .O(N__20244),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__2208 (
            .O(N__20241),
            .I(N__20238));
    LocalMux I__2207 (
            .O(N__20238),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__2206 (
            .O(N__20235),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ));
    InMux I__2205 (
            .O(N__20232),
            .I(N__20229));
    LocalMux I__2204 (
            .O(N__20229),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2203 (
            .O(N__20226),
            .I(N__20223));
    LocalMux I__2202 (
            .O(N__20223),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9 ));
    InMux I__2201 (
            .O(N__20220),
            .I(N__20215));
    InMux I__2200 (
            .O(N__20219),
            .I(N__20212));
    InMux I__2199 (
            .O(N__20218),
            .I(N__20209));
    LocalMux I__2198 (
            .O(N__20215),
            .I(N__20206));
    LocalMux I__2197 (
            .O(N__20212),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__2196 (
            .O(N__20209),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    Odrv4 I__2195 (
            .O(N__20206),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    CascadeMux I__2194 (
            .O(N__20199),
            .I(N__20196));
    InMux I__2193 (
            .O(N__20196),
            .I(N__20193));
    LocalMux I__2192 (
            .O(N__20193),
            .I(N__20190));
    Span4Mux_s3_h I__2191 (
            .O(N__20190),
            .I(N__20187));
    Odrv4 I__2190 (
            .O(N__20187),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    InMux I__2189 (
            .O(N__20184),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__2188 (
            .O(N__20181),
            .I(N__20178));
    LocalMux I__2187 (
            .O(N__20178),
            .I(N__20174));
    InMux I__2186 (
            .O(N__20177),
            .I(N__20171));
    Span4Mux_v I__2185 (
            .O(N__20174),
            .I(N__20168));
    LocalMux I__2184 (
            .O(N__20171),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    Odrv4 I__2183 (
            .O(N__20168),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    InMux I__2182 (
            .O(N__20163),
            .I(N__20160));
    LocalMux I__2181 (
            .O(N__20160),
            .I(N__20157));
    Span4Mux_s3_h I__2180 (
            .O(N__20157),
            .I(N__20154));
    Odrv4 I__2179 (
            .O(N__20154),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__2178 (
            .O(N__20151),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__2177 (
            .O(N__20148),
            .I(N__20141));
    InMux I__2176 (
            .O(N__20147),
            .I(N__20141));
    InMux I__2175 (
            .O(N__20146),
            .I(N__20138));
    LocalMux I__2174 (
            .O(N__20141),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__2173 (
            .O(N__20138),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__2172 (
            .O(N__20133),
            .I(N__20130));
    LocalMux I__2171 (
            .O(N__20130),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    InMux I__2170 (
            .O(N__20127),
            .I(bfn_3_13_0_));
    CascadeMux I__2169 (
            .O(N__20124),
            .I(N__20121));
    InMux I__2168 (
            .O(N__20121),
            .I(N__20118));
    LocalMux I__2167 (
            .O(N__20118),
            .I(N__20113));
    InMux I__2166 (
            .O(N__20117),
            .I(N__20110));
    InMux I__2165 (
            .O(N__20116),
            .I(N__20107));
    Span4Mux_v I__2164 (
            .O(N__20113),
            .I(N__20104));
    LocalMux I__2163 (
            .O(N__20110),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__2162 (
            .O(N__20107),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    Odrv4 I__2161 (
            .O(N__20104),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__2160 (
            .O(N__20097),
            .I(N__20094));
    LocalMux I__2159 (
            .O(N__20094),
            .I(N__20091));
    Span4Mux_h I__2158 (
            .O(N__20091),
            .I(N__20088));
    Odrv4 I__2157 (
            .O(N__20088),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    InMux I__2156 (
            .O(N__20085),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__2155 (
            .O(N__20082),
            .I(N__20078));
    CascadeMux I__2154 (
            .O(N__20081),
            .I(N__20074));
    LocalMux I__2153 (
            .O(N__20078),
            .I(N__20071));
    InMux I__2152 (
            .O(N__20077),
            .I(N__20068));
    InMux I__2151 (
            .O(N__20074),
            .I(N__20065));
    Span4Mux_v I__2150 (
            .O(N__20071),
            .I(N__20062));
    LocalMux I__2149 (
            .O(N__20068),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    LocalMux I__2148 (
            .O(N__20065),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    Odrv4 I__2147 (
            .O(N__20062),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__2146 (
            .O(N__20055),
            .I(N__20052));
    LocalMux I__2145 (
            .O(N__20052),
            .I(N__20049));
    Odrv4 I__2144 (
            .O(N__20049),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    InMux I__2143 (
            .O(N__20046),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__2142 (
            .O(N__20043),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__2141 (
            .O(N__20040),
            .I(N__20037));
    LocalMux I__2140 (
            .O(N__20037),
            .I(N__20034));
    Odrv12 I__2139 (
            .O(N__20034),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    InMux I__2138 (
            .O(N__20031),
            .I(N__20028));
    LocalMux I__2137 (
            .O(N__20028),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__2136 (
            .O(N__20025),
            .I(N__20022));
    LocalMux I__2135 (
            .O(N__20022),
            .I(N__20019));
    Span4Mux_v I__2134 (
            .O(N__20019),
            .I(N__20016));
    Odrv4 I__2133 (
            .O(N__20016),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__2132 (
            .O(N__20013),
            .I(N__20010));
    LocalMux I__2131 (
            .O(N__20010),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    InMux I__2130 (
            .O(N__20007),
            .I(N__20004));
    LocalMux I__2129 (
            .O(N__20004),
            .I(N__20001));
    Span4Mux_h I__2128 (
            .O(N__20001),
            .I(N__19998));
    Odrv4 I__2127 (
            .O(N__19998),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__2126 (
            .O(N__19995),
            .I(N__19992));
    LocalMux I__2125 (
            .O(N__19992),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__2124 (
            .O(N__19989),
            .I(N__19986));
    LocalMux I__2123 (
            .O(N__19986),
            .I(N__19983));
    Span4Mux_h I__2122 (
            .O(N__19983),
            .I(N__19980));
    Odrv4 I__2121 (
            .O(N__19980),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__2120 (
            .O(N__19977),
            .I(N__19974));
    LocalMux I__2119 (
            .O(N__19974),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__2118 (
            .O(N__19971),
            .I(N__19968));
    LocalMux I__2117 (
            .O(N__19968),
            .I(N__19965));
    Span4Mux_h I__2116 (
            .O(N__19965),
            .I(N__19962));
    Odrv4 I__2115 (
            .O(N__19962),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__2114 (
            .O(N__19959),
            .I(N__19956));
    LocalMux I__2113 (
            .O(N__19956),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__2112 (
            .O(N__19953),
            .I(N__19949));
    InMux I__2111 (
            .O(N__19952),
            .I(N__19945));
    LocalMux I__2110 (
            .O(N__19949),
            .I(N__19942));
    InMux I__2109 (
            .O(N__19948),
            .I(N__19939));
    LocalMux I__2108 (
            .O(N__19945),
            .I(N__19936));
    Span4Mux_v I__2107 (
            .O(N__19942),
            .I(N__19933));
    LocalMux I__2106 (
            .O(N__19939),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    Odrv4 I__2105 (
            .O(N__19936),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    Odrv4 I__2104 (
            .O(N__19933),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    CascadeMux I__2103 (
            .O(N__19926),
            .I(N__19923));
    InMux I__2102 (
            .O(N__19923),
            .I(N__19920));
    LocalMux I__2101 (
            .O(N__19920),
            .I(N__19917));
    Odrv4 I__2100 (
            .O(N__19917),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    InMux I__2099 (
            .O(N__19914),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    CascadeMux I__2098 (
            .O(N__19911),
            .I(N__19906));
    CascadeMux I__2097 (
            .O(N__19910),
            .I(N__19901));
    InMux I__2096 (
            .O(N__19909),
            .I(N__19897));
    InMux I__2095 (
            .O(N__19906),
            .I(N__19894));
    InMux I__2094 (
            .O(N__19905),
            .I(N__19887));
    InMux I__2093 (
            .O(N__19904),
            .I(N__19880));
    InMux I__2092 (
            .O(N__19901),
            .I(N__19880));
    InMux I__2091 (
            .O(N__19900),
            .I(N__19880));
    LocalMux I__2090 (
            .O(N__19897),
            .I(N__19875));
    LocalMux I__2089 (
            .O(N__19894),
            .I(N__19875));
    InMux I__2088 (
            .O(N__19893),
            .I(N__19866));
    InMux I__2087 (
            .O(N__19892),
            .I(N__19866));
    InMux I__2086 (
            .O(N__19891),
            .I(N__19866));
    InMux I__2085 (
            .O(N__19890),
            .I(N__19866));
    LocalMux I__2084 (
            .O(N__19887),
            .I(N__19860));
    LocalMux I__2083 (
            .O(N__19880),
            .I(N__19860));
    Span4Mux_h I__2082 (
            .O(N__19875),
            .I(N__19855));
    LocalMux I__2081 (
            .O(N__19866),
            .I(N__19855));
    InMux I__2080 (
            .O(N__19865),
            .I(N__19852));
    Odrv4 I__2079 (
            .O(N__19860),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2078 (
            .O(N__19855),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2077 (
            .O(N__19852),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    InMux I__2076 (
            .O(N__19845),
            .I(N__19842));
    LocalMux I__2075 (
            .O(N__19842),
            .I(N__19838));
    InMux I__2074 (
            .O(N__19841),
            .I(N__19835));
    Span4Mux_h I__2073 (
            .O(N__19838),
            .I(N__19830));
    LocalMux I__2072 (
            .O(N__19835),
            .I(N__19830));
    Odrv4 I__2071 (
            .O(N__19830),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__2070 (
            .O(N__19827),
            .I(N__19824));
    LocalMux I__2069 (
            .O(N__19824),
            .I(N__19821));
    Odrv12 I__2068 (
            .O(N__19821),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__2067 (
            .O(N__19818),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    InMux I__2066 (
            .O(N__19815),
            .I(N__19812));
    LocalMux I__2065 (
            .O(N__19812),
            .I(N__19807));
    InMux I__2064 (
            .O(N__19811),
            .I(N__19804));
    InMux I__2063 (
            .O(N__19810),
            .I(N__19801));
    Span4Mux_v I__2062 (
            .O(N__19807),
            .I(N__19798));
    LocalMux I__2061 (
            .O(N__19804),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__2060 (
            .O(N__19801),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    Odrv4 I__2059 (
            .O(N__19798),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    CascadeMux I__2058 (
            .O(N__19791),
            .I(N__19788));
    InMux I__2057 (
            .O(N__19788),
            .I(N__19785));
    LocalMux I__2056 (
            .O(N__19785),
            .I(N__19782));
    Odrv4 I__2055 (
            .O(N__19782),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    InMux I__2054 (
            .O(N__19779),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    InMux I__2053 (
            .O(N__19776),
            .I(N__19772));
    InMux I__2052 (
            .O(N__19775),
            .I(N__19769));
    LocalMux I__2051 (
            .O(N__19772),
            .I(N__19766));
    LocalMux I__2050 (
            .O(N__19769),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    Odrv4 I__2049 (
            .O(N__19766),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    InMux I__2048 (
            .O(N__19761),
            .I(N__19758));
    LocalMux I__2047 (
            .O(N__19758),
            .I(N__19755));
    Span4Mux_v I__2046 (
            .O(N__19755),
            .I(N__19752));
    Odrv4 I__2045 (
            .O(N__19752),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    InMux I__2044 (
            .O(N__19749),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__2043 (
            .O(N__19746),
            .I(N__19743));
    LocalMux I__2042 (
            .O(N__19743),
            .I(N__19740));
    Span4Mux_h I__2041 (
            .O(N__19740),
            .I(N__19736));
    InMux I__2040 (
            .O(N__19739),
            .I(N__19733));
    Odrv4 I__2039 (
            .O(N__19736),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    LocalMux I__2038 (
            .O(N__19733),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    CascadeMux I__2037 (
            .O(N__19728),
            .I(N__19725));
    InMux I__2036 (
            .O(N__19725),
            .I(N__19722));
    LocalMux I__2035 (
            .O(N__19722),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    InMux I__2034 (
            .O(N__19719),
            .I(N__19716));
    LocalMux I__2033 (
            .O(N__19716),
            .I(N__19713));
    Span4Mux_h I__2032 (
            .O(N__19713),
            .I(N__19710));
    Odrv4 I__2031 (
            .O(N__19710),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__2030 (
            .O(N__19707),
            .I(N__19704));
    LocalMux I__2029 (
            .O(N__19704),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__2028 (
            .O(N__19701),
            .I(N__19698));
    LocalMux I__2027 (
            .O(N__19698),
            .I(N__19695));
    Span4Mux_v I__2026 (
            .O(N__19695),
            .I(N__19692));
    Odrv4 I__2025 (
            .O(N__19692),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__2024 (
            .O(N__19689),
            .I(N__19686));
    LocalMux I__2023 (
            .O(N__19686),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__2022 (
            .O(N__19683),
            .I(N__19680));
    LocalMux I__2021 (
            .O(N__19680),
            .I(N__19677));
    Span4Mux_h I__2020 (
            .O(N__19677),
            .I(N__19674));
    Odrv4 I__2019 (
            .O(N__19674),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__2018 (
            .O(N__19671),
            .I(N__19668));
    LocalMux I__2017 (
            .O(N__19668),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__2016 (
            .O(N__19665),
            .I(N__19662));
    LocalMux I__2015 (
            .O(N__19662),
            .I(N__19659));
    Span4Mux_h I__2014 (
            .O(N__19659),
            .I(N__19656));
    Odrv4 I__2013 (
            .O(N__19656),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__2012 (
            .O(N__19653),
            .I(N__19650));
    LocalMux I__2011 (
            .O(N__19650),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__2010 (
            .O(N__19647),
            .I(N__19644));
    LocalMux I__2009 (
            .O(N__19644),
            .I(N__19641));
    Span4Mux_v I__2008 (
            .O(N__19641),
            .I(N__19638));
    Span4Mux_h I__2007 (
            .O(N__19638),
            .I(N__19635));
    Odrv4 I__2006 (
            .O(N__19635),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__2005 (
            .O(N__19632),
            .I(N__19629));
    LocalMux I__2004 (
            .O(N__19629),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__2003 (
            .O(N__19626),
            .I(N__19623));
    LocalMux I__2002 (
            .O(N__19623),
            .I(N__19620));
    Span12Mux_v I__2001 (
            .O(N__19620),
            .I(N__19617));
    Odrv12 I__2000 (
            .O(N__19617),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1999 (
            .O(N__19614),
            .I(N__19611));
    LocalMux I__1998 (
            .O(N__19611),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__1997 (
            .O(N__19608),
            .I(N__19605));
    LocalMux I__1996 (
            .O(N__19605),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__1995 (
            .O(N__19602),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__1994 (
            .O(N__19599),
            .I(N__19596));
    LocalMux I__1993 (
            .O(N__19596),
            .I(N__19593));
    Span4Mux_h I__1992 (
            .O(N__19593),
            .I(N__19590));
    Odrv4 I__1991 (
            .O(N__19590),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__1990 (
            .O(N__19587),
            .I(N__19584));
    LocalMux I__1989 (
            .O(N__19584),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__1988 (
            .O(N__19581),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__1987 (
            .O(N__19578),
            .I(N__19575));
    LocalMux I__1986 (
            .O(N__19575),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    InMux I__1985 (
            .O(N__19572),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    InMux I__1984 (
            .O(N__19569),
            .I(bfn_3_9_0_));
    CascadeMux I__1983 (
            .O(N__19566),
            .I(N__19563));
    InMux I__1982 (
            .O(N__19563),
            .I(N__19560));
    LocalMux I__1981 (
            .O(N__19560),
            .I(N__19557));
    Span4Mux_v I__1980 (
            .O(N__19557),
            .I(N__19554));
    Odrv4 I__1979 (
            .O(N__19554),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__1978 (
            .O(N__19551),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    InMux I__1977 (
            .O(N__19548),
            .I(N__19545));
    LocalMux I__1976 (
            .O(N__19545),
            .I(N__19541));
    InMux I__1975 (
            .O(N__19544),
            .I(N__19538));
    Odrv4 I__1974 (
            .O(N__19541),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    LocalMux I__1973 (
            .O(N__19538),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    InMux I__1972 (
            .O(N__19533),
            .I(N__19530));
    LocalMux I__1971 (
            .O(N__19530),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    InMux I__1970 (
            .O(N__19527),
            .I(N__19523));
    InMux I__1969 (
            .O(N__19526),
            .I(N__19520));
    LocalMux I__1968 (
            .O(N__19523),
            .I(N__19517));
    LocalMux I__1967 (
            .O(N__19520),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    Odrv4 I__1966 (
            .O(N__19517),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__1965 (
            .O(N__19512),
            .I(N__19509));
    LocalMux I__1964 (
            .O(N__19509),
            .I(N__19505));
    InMux I__1963 (
            .O(N__19508),
            .I(N__19502));
    Odrv4 I__1962 (
            .O(N__19505),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    LocalMux I__1961 (
            .O(N__19502),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    InMux I__1960 (
            .O(N__19497),
            .I(N__19494));
    LocalMux I__1959 (
            .O(N__19494),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__1958 (
            .O(N__19491),
            .I(N__19488));
    LocalMux I__1957 (
            .O(N__19488),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__1956 (
            .O(N__19485),
            .I(N__19482));
    LocalMux I__1955 (
            .O(N__19482),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    InMux I__1954 (
            .O(N__19479),
            .I(N__19476));
    LocalMux I__1953 (
            .O(N__19476),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__1952 (
            .O(N__19473),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__1951 (
            .O(N__19470),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    CascadeMux I__1950 (
            .O(N__19467),
            .I(N__19464));
    InMux I__1949 (
            .O(N__19464),
            .I(N__19461));
    LocalMux I__1948 (
            .O(N__19461),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    InMux I__1947 (
            .O(N__19458),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__1946 (
            .O(N__19455),
            .I(N__19452));
    LocalMux I__1945 (
            .O(N__19452),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    InMux I__1944 (
            .O(N__19449),
            .I(N__19446));
    LocalMux I__1943 (
            .O(N__19446),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__1942 (
            .O(N__19443),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__1941 (
            .O(N__19440),
            .I(N__19437));
    LocalMux I__1940 (
            .O(N__19437),
            .I(\current_shift_inst.PI_CTRL.N_98 ));
    InMux I__1939 (
            .O(N__19434),
            .I(N__19424));
    InMux I__1938 (
            .O(N__19433),
            .I(N__19424));
    InMux I__1937 (
            .O(N__19432),
            .I(N__19424));
    InMux I__1936 (
            .O(N__19431),
            .I(N__19421));
    LocalMux I__1935 (
            .O(N__19424),
            .I(N__19415));
    LocalMux I__1934 (
            .O(N__19421),
            .I(N__19415));
    InMux I__1933 (
            .O(N__19420),
            .I(N__19412));
    Span4Mux_v I__1932 (
            .O(N__19415),
            .I(N__19409));
    LocalMux I__1931 (
            .O(N__19412),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    Odrv4 I__1930 (
            .O(N__19409),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    CascadeMux I__1929 (
            .O(N__19404),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_ ));
    InMux I__1928 (
            .O(N__19401),
            .I(N__19392));
    InMux I__1927 (
            .O(N__19400),
            .I(N__19383));
    InMux I__1926 (
            .O(N__19399),
            .I(N__19383));
    InMux I__1925 (
            .O(N__19398),
            .I(N__19383));
    InMux I__1924 (
            .O(N__19397),
            .I(N__19383));
    InMux I__1923 (
            .O(N__19396),
            .I(N__19377));
    InMux I__1922 (
            .O(N__19395),
            .I(N__19377));
    LocalMux I__1921 (
            .O(N__19392),
            .I(N__19371));
    LocalMux I__1920 (
            .O(N__19383),
            .I(N__19371));
    InMux I__1919 (
            .O(N__19382),
            .I(N__19368));
    LocalMux I__1918 (
            .O(N__19377),
            .I(N__19365));
    InMux I__1917 (
            .O(N__19376),
            .I(N__19362));
    Odrv4 I__1916 (
            .O(N__19371),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    LocalMux I__1915 (
            .O(N__19368),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    Odrv12 I__1914 (
            .O(N__19365),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    LocalMux I__1913 (
            .O(N__19362),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    CascadeMux I__1912 (
            .O(N__19353),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ));
    InMux I__1911 (
            .O(N__19350),
            .I(N__19346));
    InMux I__1910 (
            .O(N__19349),
            .I(N__19343));
    LocalMux I__1909 (
            .O(N__19346),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__1908 (
            .O(N__19343),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__1907 (
            .O(N__19338),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ));
    InMux I__1906 (
            .O(N__19335),
            .I(N__19332));
    LocalMux I__1905 (
            .O(N__19332),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__1904 (
            .O(N__19329),
            .I(N__19326));
    LocalMux I__1903 (
            .O(N__19326),
            .I(N__19323));
    Odrv4 I__1902 (
            .O(N__19323),
            .I(un7_start_stop_0_a3));
    InMux I__1901 (
            .O(N__19320),
            .I(N__19317));
    LocalMux I__1900 (
            .O(N__19317),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__1899 (
            .O(N__19314),
            .I(N__19311));
    LocalMux I__1898 (
            .O(N__19311),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1897 (
            .O(N__19308),
            .I(bfn_2_12_0_));
    CascadeMux I__1896 (
            .O(N__19305),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ));
    InMux I__1895 (
            .O(N__19302),
            .I(N__19298));
    InMux I__1894 (
            .O(N__19301),
            .I(N__19295));
    LocalMux I__1893 (
            .O(N__19298),
            .I(N__19292));
    LocalMux I__1892 (
            .O(N__19295),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    Odrv12 I__1891 (
            .O(N__19292),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    InMux I__1890 (
            .O(N__19287),
            .I(N__19281));
    InMux I__1889 (
            .O(N__19286),
            .I(N__19281));
    LocalMux I__1888 (
            .O(N__19281),
            .I(N__19278));
    Odrv4 I__1887 (
            .O(N__19278),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    CascadeMux I__1886 (
            .O(N__19275),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__1885 (
            .O(N__19272),
            .I(N__19269));
    LocalMux I__1884 (
            .O(N__19269),
            .I(N__19265));
    InMux I__1883 (
            .O(N__19268),
            .I(N__19262));
    Odrv12 I__1882 (
            .O(N__19265),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__1881 (
            .O(N__19262),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__1880 (
            .O(N__19257),
            .I(\current_shift_inst.PI_CTRL.N_31_cascade_ ));
    InMux I__1879 (
            .O(N__19254),
            .I(N__19251));
    LocalMux I__1878 (
            .O(N__19251),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    InMux I__1877 (
            .O(N__19248),
            .I(N__19245));
    LocalMux I__1876 (
            .O(N__19245),
            .I(N__19242));
    Span4Mux_h I__1875 (
            .O(N__19242),
            .I(N__19239));
    Odrv4 I__1874 (
            .O(N__19239),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    CascadeMux I__1873 (
            .O(N__19236),
            .I(N__19233));
    InMux I__1872 (
            .O(N__19233),
            .I(N__19230));
    LocalMux I__1871 (
            .O(N__19230),
            .I(N__19227));
    Span4Mux_h I__1870 (
            .O(N__19227),
            .I(N__19224));
    Span4Mux_v I__1869 (
            .O(N__19224),
            .I(N__19221));
    Odrv4 I__1868 (
            .O(N__19221),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    InMux I__1867 (
            .O(N__19218),
            .I(N__19215));
    LocalMux I__1866 (
            .O(N__19215),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__1865 (
            .O(N__19212),
            .I(bfn_2_11_0_));
    InMux I__1864 (
            .O(N__19209),
            .I(N__19206));
    LocalMux I__1863 (
            .O(N__19206),
            .I(N__19203));
    Span4Mux_h I__1862 (
            .O(N__19203),
            .I(N__19200));
    Odrv4 I__1861 (
            .O(N__19200),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    CascadeMux I__1860 (
            .O(N__19197),
            .I(N__19194));
    InMux I__1859 (
            .O(N__19194),
            .I(N__19191));
    LocalMux I__1858 (
            .O(N__19191),
            .I(N__19188));
    Span4Mux_h I__1857 (
            .O(N__19188),
            .I(N__19185));
    Span4Mux_v I__1856 (
            .O(N__19185),
            .I(N__19182));
    Odrv4 I__1855 (
            .O(N__19182),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    InMux I__1854 (
            .O(N__19179),
            .I(N__19176));
    LocalMux I__1853 (
            .O(N__19176),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__1852 (
            .O(N__19173),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    CascadeMux I__1851 (
            .O(N__19170),
            .I(N__19167));
    InMux I__1850 (
            .O(N__19167),
            .I(N__19164));
    LocalMux I__1849 (
            .O(N__19164),
            .I(N__19161));
    Span4Mux_h I__1848 (
            .O(N__19161),
            .I(N__19158));
    Span4Mux_v I__1847 (
            .O(N__19158),
            .I(N__19155));
    Odrv4 I__1846 (
            .O(N__19155),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1845 (
            .O(N__19152),
            .I(N__19149));
    LocalMux I__1844 (
            .O(N__19149),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__1843 (
            .O(N__19146),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    InMux I__1842 (
            .O(N__19143),
            .I(N__19140));
    LocalMux I__1841 (
            .O(N__19140),
            .I(N__19137));
    Span4Mux_h I__1840 (
            .O(N__19137),
            .I(N__19134));
    Span4Mux_v I__1839 (
            .O(N__19134),
            .I(N__19131));
    Odrv4 I__1838 (
            .O(N__19131),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1837 (
            .O(N__19128),
            .I(N__19125));
    LocalMux I__1836 (
            .O(N__19125),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__1835 (
            .O(N__19122),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    CascadeMux I__1834 (
            .O(N__19119),
            .I(N__19116));
    InMux I__1833 (
            .O(N__19116),
            .I(N__19113));
    LocalMux I__1832 (
            .O(N__19113),
            .I(N__19110));
    Span4Mux_v I__1831 (
            .O(N__19110),
            .I(N__19107));
    Span4Mux_v I__1830 (
            .O(N__19107),
            .I(N__19104));
    Odrv4 I__1829 (
            .O(N__19104),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1828 (
            .O(N__19101),
            .I(N__19098));
    LocalMux I__1827 (
            .O(N__19098),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__1826 (
            .O(N__19095),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    InMux I__1825 (
            .O(N__19092),
            .I(N__19089));
    LocalMux I__1824 (
            .O(N__19089),
            .I(N__19086));
    Span4Mux_v I__1823 (
            .O(N__19086),
            .I(N__19083));
    Span4Mux_v I__1822 (
            .O(N__19083),
            .I(N__19080));
    Odrv4 I__1821 (
            .O(N__19080),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__1820 (
            .O(N__19077),
            .I(N__19074));
    LocalMux I__1819 (
            .O(N__19074),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__1818 (
            .O(N__19071),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    CascadeMux I__1817 (
            .O(N__19068),
            .I(N__19065));
    InMux I__1816 (
            .O(N__19065),
            .I(N__19062));
    LocalMux I__1815 (
            .O(N__19062),
            .I(N__19059));
    Span4Mux_h I__1814 (
            .O(N__19059),
            .I(N__19056));
    Span4Mux_v I__1813 (
            .O(N__19056),
            .I(N__19053));
    Odrv4 I__1812 (
            .O(N__19053),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1811 (
            .O(N__19050),
            .I(N__19047));
    LocalMux I__1810 (
            .O(N__19047),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__1809 (
            .O(N__19044),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    InMux I__1808 (
            .O(N__19041),
            .I(N__19038));
    LocalMux I__1807 (
            .O(N__19038),
            .I(N__19035));
    Span4Mux_v I__1806 (
            .O(N__19035),
            .I(N__19032));
    Odrv4 I__1805 (
            .O(N__19032),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    CascadeMux I__1804 (
            .O(N__19029),
            .I(N__19022));
    CascadeMux I__1803 (
            .O(N__19028),
            .I(N__19018));
    CascadeMux I__1802 (
            .O(N__19027),
            .I(N__19014));
    InMux I__1801 (
            .O(N__19026),
            .I(N__19010));
    InMux I__1800 (
            .O(N__19025),
            .I(N__19007));
    InMux I__1799 (
            .O(N__19022),
            .I(N__18994));
    InMux I__1798 (
            .O(N__19021),
            .I(N__18994));
    InMux I__1797 (
            .O(N__19018),
            .I(N__18994));
    InMux I__1796 (
            .O(N__19017),
            .I(N__18994));
    InMux I__1795 (
            .O(N__19014),
            .I(N__18994));
    InMux I__1794 (
            .O(N__19013),
            .I(N__18994));
    LocalMux I__1793 (
            .O(N__19010),
            .I(N__18991));
    LocalMux I__1792 (
            .O(N__19007),
            .I(N__18986));
    LocalMux I__1791 (
            .O(N__18994),
            .I(N__18986));
    Span4Mux_v I__1790 (
            .O(N__18991),
            .I(N__18983));
    Span4Mux_h I__1789 (
            .O(N__18986),
            .I(N__18980));
    Odrv4 I__1788 (
            .O(N__18983),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    Odrv4 I__1787 (
            .O(N__18980),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    InMux I__1786 (
            .O(N__18975),
            .I(N__18972));
    LocalMux I__1785 (
            .O(N__18972),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__1784 (
            .O(N__18969),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1783 (
            .O(N__18966),
            .I(N__18963));
    LocalMux I__1782 (
            .O(N__18963),
            .I(N__18960));
    Span4Mux_h I__1781 (
            .O(N__18960),
            .I(N__18957));
    Odrv4 I__1780 (
            .O(N__18957),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    CascadeMux I__1779 (
            .O(N__18954),
            .I(N__18951));
    InMux I__1778 (
            .O(N__18951),
            .I(N__18948));
    LocalMux I__1777 (
            .O(N__18948),
            .I(N__18945));
    Span4Mux_h I__1776 (
            .O(N__18945),
            .I(N__18942));
    Span4Mux_v I__1775 (
            .O(N__18942),
            .I(N__18939));
    Odrv4 I__1774 (
            .O(N__18939),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    CascadeMux I__1773 (
            .O(N__18936),
            .I(N__18933));
    InMux I__1772 (
            .O(N__18933),
            .I(N__18930));
    LocalMux I__1771 (
            .O(N__18930),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__1770 (
            .O(N__18927),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1769 (
            .O(N__18924),
            .I(N__18921));
    LocalMux I__1768 (
            .O(N__18921),
            .I(N__18918));
    Span4Mux_h I__1767 (
            .O(N__18918),
            .I(N__18915));
    Odrv4 I__1766 (
            .O(N__18915),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    CascadeMux I__1765 (
            .O(N__18912),
            .I(N__18909));
    InMux I__1764 (
            .O(N__18909),
            .I(N__18906));
    LocalMux I__1763 (
            .O(N__18906),
            .I(N__18903));
    Span4Mux_h I__1762 (
            .O(N__18903),
            .I(N__18900));
    Span4Mux_v I__1761 (
            .O(N__18900),
            .I(N__18897));
    Odrv4 I__1760 (
            .O(N__18897),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    InMux I__1759 (
            .O(N__18894),
            .I(N__18891));
    LocalMux I__1758 (
            .O(N__18891),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__1757 (
            .O(N__18888),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1756 (
            .O(N__18885),
            .I(N__18882));
    LocalMux I__1755 (
            .O(N__18882),
            .I(N__18879));
    Span4Mux_v I__1754 (
            .O(N__18879),
            .I(N__18876));
    Odrv4 I__1753 (
            .O(N__18876),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    CascadeMux I__1752 (
            .O(N__18873),
            .I(N__18870));
    InMux I__1751 (
            .O(N__18870),
            .I(N__18867));
    LocalMux I__1750 (
            .O(N__18867),
            .I(N__18864));
    Span4Mux_h I__1749 (
            .O(N__18864),
            .I(N__18861));
    Span4Mux_v I__1748 (
            .O(N__18861),
            .I(N__18858));
    Odrv4 I__1747 (
            .O(N__18858),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    InMux I__1746 (
            .O(N__18855),
            .I(N__18852));
    LocalMux I__1745 (
            .O(N__18852),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__1744 (
            .O(N__18849),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1743 (
            .O(N__18846),
            .I(N__18843));
    LocalMux I__1742 (
            .O(N__18843),
            .I(N__18840));
    Span4Mux_v I__1741 (
            .O(N__18840),
            .I(N__18837));
    Odrv4 I__1740 (
            .O(N__18837),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    CascadeMux I__1739 (
            .O(N__18834),
            .I(N__18831));
    InMux I__1738 (
            .O(N__18831),
            .I(N__18828));
    LocalMux I__1737 (
            .O(N__18828),
            .I(N__18825));
    Span4Mux_v I__1736 (
            .O(N__18825),
            .I(N__18822));
    Span4Mux_v I__1735 (
            .O(N__18822),
            .I(N__18819));
    Odrv4 I__1734 (
            .O(N__18819),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    InMux I__1733 (
            .O(N__18816),
            .I(N__18813));
    LocalMux I__1732 (
            .O(N__18813),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__1731 (
            .O(N__18810),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1730 (
            .O(N__18807),
            .I(N__18804));
    LocalMux I__1729 (
            .O(N__18804),
            .I(N__18801));
    Span4Mux_h I__1728 (
            .O(N__18801),
            .I(N__18798));
    Odrv4 I__1727 (
            .O(N__18798),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    CascadeMux I__1726 (
            .O(N__18795),
            .I(N__18792));
    InMux I__1725 (
            .O(N__18792),
            .I(N__18789));
    LocalMux I__1724 (
            .O(N__18789),
            .I(N__18786));
    Span4Mux_v I__1723 (
            .O(N__18786),
            .I(N__18783));
    Span4Mux_v I__1722 (
            .O(N__18783),
            .I(N__18780));
    Odrv4 I__1721 (
            .O(N__18780),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    InMux I__1720 (
            .O(N__18777),
            .I(N__18774));
    LocalMux I__1719 (
            .O(N__18774),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__1718 (
            .O(N__18771),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1717 (
            .O(N__18768),
            .I(N__18765));
    LocalMux I__1716 (
            .O(N__18765),
            .I(N__18762));
    Span4Mux_h I__1715 (
            .O(N__18762),
            .I(N__18759));
    Odrv4 I__1714 (
            .O(N__18759),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    CascadeMux I__1713 (
            .O(N__18756),
            .I(N__18753));
    InMux I__1712 (
            .O(N__18753),
            .I(N__18750));
    LocalMux I__1711 (
            .O(N__18750),
            .I(N__18747));
    Span4Mux_h I__1710 (
            .O(N__18747),
            .I(N__18744));
    Span4Mux_v I__1709 (
            .O(N__18744),
            .I(N__18741));
    Odrv4 I__1708 (
            .O(N__18741),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    InMux I__1707 (
            .O(N__18738),
            .I(N__18735));
    LocalMux I__1706 (
            .O(N__18735),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__1705 (
            .O(N__18732),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1704 (
            .O(N__18729),
            .I(N__18726));
    LocalMux I__1703 (
            .O(N__18726),
            .I(N__18723));
    Span4Mux_h I__1702 (
            .O(N__18723),
            .I(N__18720));
    Odrv4 I__1701 (
            .O(N__18720),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    CascadeMux I__1700 (
            .O(N__18717),
            .I(N__18714));
    InMux I__1699 (
            .O(N__18714),
            .I(N__18711));
    LocalMux I__1698 (
            .O(N__18711),
            .I(N__18708));
    Span4Mux_h I__1697 (
            .O(N__18708),
            .I(N__18705));
    Span4Mux_v I__1696 (
            .O(N__18705),
            .I(N__18702));
    Odrv4 I__1695 (
            .O(N__18702),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    InMux I__1694 (
            .O(N__18699),
            .I(N__18696));
    LocalMux I__1693 (
            .O(N__18696),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__1692 (
            .O(N__18693),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1691 (
            .O(N__18690),
            .I(N__18684));
    InMux I__1690 (
            .O(N__18689),
            .I(N__18684));
    LocalMux I__1689 (
            .O(N__18684),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    CascadeMux I__1688 (
            .O(N__18681),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ));
    InMux I__1687 (
            .O(N__18678),
            .I(N__18675));
    LocalMux I__1686 (
            .O(N__18675),
            .I(N__18672));
    Span4Mux_v I__1685 (
            .O(N__18672),
            .I(N__18668));
    InMux I__1684 (
            .O(N__18671),
            .I(N__18665));
    Odrv4 I__1683 (
            .O(N__18668),
            .I(\pwm_generator_inst.O_10 ));
    LocalMux I__1682 (
            .O(N__18665),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1681 (
            .O(N__18660),
            .I(N__18654));
    InMux I__1680 (
            .O(N__18659),
            .I(N__18654));
    LocalMux I__1679 (
            .O(N__18654),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    CascadeMux I__1678 (
            .O(N__18651),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_ ));
    InMux I__1677 (
            .O(N__18648),
            .I(N__18645));
    LocalMux I__1676 (
            .O(N__18645),
            .I(N__18642));
    Span4Mux_h I__1675 (
            .O(N__18642),
            .I(N__18639));
    Span4Mux_v I__1674 (
            .O(N__18639),
            .I(N__18636));
    Odrv4 I__1673 (
            .O(N__18636),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1672 (
            .O(N__18633),
            .I(N__18630));
    InMux I__1671 (
            .O(N__18630),
            .I(N__18627));
    LocalMux I__1670 (
            .O(N__18627),
            .I(N__18624));
    Span4Mux_h I__1669 (
            .O(N__18624),
            .I(N__18621));
    Odrv4 I__1668 (
            .O(N__18621),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1667 (
            .O(N__18618),
            .I(N__18615));
    LocalMux I__1666 (
            .O(N__18615),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    InMux I__1665 (
            .O(N__18612),
            .I(N__18606));
    InMux I__1664 (
            .O(N__18611),
            .I(N__18606));
    LocalMux I__1663 (
            .O(N__18606),
            .I(N__18602));
    InMux I__1662 (
            .O(N__18605),
            .I(N__18599));
    Odrv12 I__1661 (
            .O(N__18602),
            .I(pwm_duty_input_9));
    LocalMux I__1660 (
            .O(N__18599),
            .I(pwm_duty_input_9));
    CascadeMux I__1659 (
            .O(N__18594),
            .I(N__18590));
    InMux I__1658 (
            .O(N__18593),
            .I(N__18585));
    InMux I__1657 (
            .O(N__18590),
            .I(N__18585));
    LocalMux I__1656 (
            .O(N__18585),
            .I(N__18581));
    InMux I__1655 (
            .O(N__18584),
            .I(N__18578));
    Odrv12 I__1654 (
            .O(N__18581),
            .I(pwm_duty_input_8));
    LocalMux I__1653 (
            .O(N__18578),
            .I(pwm_duty_input_8));
    InMux I__1652 (
            .O(N__18573),
            .I(N__18570));
    LocalMux I__1651 (
            .O(N__18570),
            .I(N_22_i_i));
    InMux I__1650 (
            .O(N__18567),
            .I(N__18564));
    LocalMux I__1649 (
            .O(N__18564),
            .I(\current_shift_inst.PI_CTRL.m14_2 ));
    InMux I__1648 (
            .O(N__18561),
            .I(N__18550));
    InMux I__1647 (
            .O(N__18560),
            .I(N__18550));
    InMux I__1646 (
            .O(N__18559),
            .I(N__18547));
    InMux I__1645 (
            .O(N__18558),
            .I(N__18540));
    InMux I__1644 (
            .O(N__18557),
            .I(N__18540));
    InMux I__1643 (
            .O(N__18556),
            .I(N__18540));
    CascadeMux I__1642 (
            .O(N__18555),
            .I(N__18537));
    LocalMux I__1641 (
            .O(N__18550),
            .I(N__18517));
    LocalMux I__1640 (
            .O(N__18547),
            .I(N__18512));
    LocalMux I__1639 (
            .O(N__18540),
            .I(N__18512));
    InMux I__1638 (
            .O(N__18537),
            .I(N__18509));
    InMux I__1637 (
            .O(N__18536),
            .I(N__18506));
    InMux I__1636 (
            .O(N__18535),
            .I(N__18503));
    InMux I__1635 (
            .O(N__18534),
            .I(N__18486));
    InMux I__1634 (
            .O(N__18533),
            .I(N__18486));
    InMux I__1633 (
            .O(N__18532),
            .I(N__18486));
    InMux I__1632 (
            .O(N__18531),
            .I(N__18486));
    InMux I__1631 (
            .O(N__18530),
            .I(N__18486));
    InMux I__1630 (
            .O(N__18529),
            .I(N__18486));
    InMux I__1629 (
            .O(N__18528),
            .I(N__18486));
    InMux I__1628 (
            .O(N__18527),
            .I(N__18486));
    InMux I__1627 (
            .O(N__18526),
            .I(N__18471));
    InMux I__1626 (
            .O(N__18525),
            .I(N__18471));
    InMux I__1625 (
            .O(N__18524),
            .I(N__18471));
    InMux I__1624 (
            .O(N__18523),
            .I(N__18471));
    InMux I__1623 (
            .O(N__18522),
            .I(N__18471));
    InMux I__1622 (
            .O(N__18521),
            .I(N__18471));
    InMux I__1621 (
            .O(N__18520),
            .I(N__18471));
    Span4Mux_v I__1620 (
            .O(N__18517),
            .I(N__18466));
    Span4Mux_v I__1619 (
            .O(N__18512),
            .I(N__18466));
    LocalMux I__1618 (
            .O(N__18509),
            .I(pwm_duty_input_10));
    LocalMux I__1617 (
            .O(N__18506),
            .I(pwm_duty_input_10));
    LocalMux I__1616 (
            .O(N__18503),
            .I(pwm_duty_input_10));
    LocalMux I__1615 (
            .O(N__18486),
            .I(pwm_duty_input_10));
    LocalMux I__1614 (
            .O(N__18471),
            .I(pwm_duty_input_10));
    Odrv4 I__1613 (
            .O(N__18466),
            .I(pwm_duty_input_10));
    InMux I__1612 (
            .O(N__18453),
            .I(N__18448));
    CascadeMux I__1611 (
            .O(N__18452),
            .I(N__18445));
    InMux I__1610 (
            .O(N__18451),
            .I(N__18442));
    LocalMux I__1609 (
            .O(N__18448),
            .I(N__18439));
    InMux I__1608 (
            .O(N__18445),
            .I(N__18436));
    LocalMux I__1607 (
            .O(N__18442),
            .I(N__18433));
    Span4Mux_v I__1606 (
            .O(N__18439),
            .I(N__18430));
    LocalMux I__1605 (
            .O(N__18436),
            .I(N__18427));
    Span4Mux_s1_h I__1604 (
            .O(N__18433),
            .I(N__18424));
    Odrv4 I__1603 (
            .O(N__18430),
            .I(pwm_duty_input_4));
    Odrv12 I__1602 (
            .O(N__18427),
            .I(pwm_duty_input_4));
    Odrv4 I__1601 (
            .O(N__18424),
            .I(pwm_duty_input_4));
    InMux I__1600 (
            .O(N__18417),
            .I(N__18414));
    LocalMux I__1599 (
            .O(N__18414),
            .I(N__18410));
    InMux I__1598 (
            .O(N__18413),
            .I(N__18407));
    Span4Mux_v I__1597 (
            .O(N__18410),
            .I(N__18404));
    LocalMux I__1596 (
            .O(N__18407),
            .I(pwm_duty_input_1));
    Odrv4 I__1595 (
            .O(N__18404),
            .I(pwm_duty_input_1));
    InMux I__1594 (
            .O(N__18399),
            .I(N__18396));
    LocalMux I__1593 (
            .O(N__18396),
            .I(N__18392));
    InMux I__1592 (
            .O(N__18395),
            .I(N__18389));
    Span4Mux_v I__1591 (
            .O(N__18392),
            .I(N__18386));
    LocalMux I__1590 (
            .O(N__18389),
            .I(pwm_duty_input_2));
    Odrv4 I__1589 (
            .O(N__18386),
            .I(pwm_duty_input_2));
    CascadeMux I__1588 (
            .O(N__18381),
            .I(N__18377));
    InMux I__1587 (
            .O(N__18380),
            .I(N__18374));
    InMux I__1586 (
            .O(N__18377),
            .I(N__18371));
    LocalMux I__1585 (
            .O(N__18374),
            .I(N__18368));
    LocalMux I__1584 (
            .O(N__18371),
            .I(N__18363));
    Span4Mux_v I__1583 (
            .O(N__18368),
            .I(N__18363));
    Odrv4 I__1582 (
            .O(N__18363),
            .I(pwm_duty_input_0));
    InMux I__1581 (
            .O(N__18360),
            .I(N__18356));
    InMux I__1580 (
            .O(N__18359),
            .I(N__18353));
    LocalMux I__1579 (
            .O(N__18356),
            .I(N__18350));
    LocalMux I__1578 (
            .O(N__18353),
            .I(N__18346));
    Span4Mux_h I__1577 (
            .O(N__18350),
            .I(N__18343));
    InMux I__1576 (
            .O(N__18349),
            .I(N__18340));
    Odrv12 I__1575 (
            .O(N__18346),
            .I(pwm_duty_input_3));
    Odrv4 I__1574 (
            .O(N__18343),
            .I(pwm_duty_input_3));
    LocalMux I__1573 (
            .O(N__18340),
            .I(pwm_duty_input_3));
    InMux I__1572 (
            .O(N__18333),
            .I(N__18330));
    LocalMux I__1571 (
            .O(N__18330),
            .I(\current_shift_inst.PI_CTRL.N_19 ));
    InMux I__1570 (
            .O(N__18327),
            .I(N__18318));
    InMux I__1569 (
            .O(N__18326),
            .I(N__18318));
    InMux I__1568 (
            .O(N__18325),
            .I(N__18318));
    LocalMux I__1567 (
            .O(N__18318),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__1566 (
            .O(N__18315),
            .I(N__18306));
    InMux I__1565 (
            .O(N__18314),
            .I(N__18306));
    InMux I__1564 (
            .O(N__18313),
            .I(N__18306));
    LocalMux I__1563 (
            .O(N__18306),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1562 (
            .O(N__18303),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__1561 (
            .O(N__18300),
            .I(N__18297));
    LocalMux I__1560 (
            .O(N__18297),
            .I(N__18294));
    Span4Mux_v I__1559 (
            .O(N__18294),
            .I(N__18290));
    InMux I__1558 (
            .O(N__18293),
            .I(N__18287));
    Odrv4 I__1557 (
            .O(N__18290),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    LocalMux I__1556 (
            .O(N__18287),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    CascadeMux I__1555 (
            .O(N__18282),
            .I(N__18279));
    InMux I__1554 (
            .O(N__18279),
            .I(N__18276));
    LocalMux I__1553 (
            .O(N__18276),
            .I(N__18273));
    Span4Mux_v I__1552 (
            .O(N__18273),
            .I(N__18270));
    Odrv4 I__1551 (
            .O(N__18270),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    InMux I__1550 (
            .O(N__18267),
            .I(N__18261));
    InMux I__1549 (
            .O(N__18266),
            .I(N__18261));
    LocalMux I__1548 (
            .O(N__18261),
            .I(N__18257));
    InMux I__1547 (
            .O(N__18260),
            .I(N__18254));
    Odrv12 I__1546 (
            .O(N__18257),
            .I(pwm_duty_input_7));
    LocalMux I__1545 (
            .O(N__18254),
            .I(pwm_duty_input_7));
    InMux I__1544 (
            .O(N__18249),
            .I(N__18243));
    InMux I__1543 (
            .O(N__18248),
            .I(N__18243));
    LocalMux I__1542 (
            .O(N__18243),
            .I(N__18239));
    InMux I__1541 (
            .O(N__18242),
            .I(N__18236));
    Odrv12 I__1540 (
            .O(N__18239),
            .I(pwm_duty_input_5));
    LocalMux I__1539 (
            .O(N__18236),
            .I(pwm_duty_input_5));
    InMux I__1538 (
            .O(N__18231),
            .I(bfn_1_10_0_));
    InMux I__1537 (
            .O(N__18228),
            .I(N__18225));
    LocalMux I__1536 (
            .O(N__18225),
            .I(N__18222));
    Odrv4 I__1535 (
            .O(N__18222),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1534 (
            .O(N__18219),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    InMux I__1533 (
            .O(N__18216),
            .I(N__18213));
    LocalMux I__1532 (
            .O(N__18213),
            .I(N__18210));
    Odrv4 I__1531 (
            .O(N__18210),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1530 (
            .O(N__18207),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1529 (
            .O(N__18204),
            .I(N__18201));
    LocalMux I__1528 (
            .O(N__18201),
            .I(N__18198));
    Odrv4 I__1527 (
            .O(N__18198),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1526 (
            .O(N__18195),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    InMux I__1525 (
            .O(N__18192),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    InMux I__1524 (
            .O(N__18189),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__1523 (
            .O(N__18186),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    InMux I__1522 (
            .O(N__18183),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    CascadeMux I__1521 (
            .O(N__18180),
            .I(\current_shift_inst.PI_CTRL.m7_2_cascade_ ));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_6 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_14 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_22 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_30 ),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(un5_counter_cry_8),
            .carryinitout(bfn_4_6_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_8 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_16 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_24 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_3_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_11_0_));
    defparam IN_MUX_bfv_3_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_12_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_3_12_0_));
    defparam IN_MUX_bfv_3_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_13_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_3_13_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_3_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_8_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_18_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_7_0_));
    defparam IN_MUX_bfv_18_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_18_8_0_));
    defparam IN_MUX_bfv_18_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_18_9_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\current_shift_inst.z_cry_7 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\current_shift_inst.z_cry_15 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\current_shift_inst.z_cry_23 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_8 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_16 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_24 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_7 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_15 ),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_7_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_22_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_23 ),
            .carryinitout(bfn_7_22_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_15 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_23 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryinitout(bfn_5_13_0_));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__33852),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_335_i_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__29022),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_187_i_g ));
    ICE_GB \current_shift_inst.timer_phase.running_RNIC90O_0  (
            .USERSIGNALTOGLOBALBUFFER(N__32373),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_phase.N_188_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__27531),
            .CLKHFEN(N__27535),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__27556),
            .RGB2PWM(N__18573),
            .RGB1(rgb_g),
            .CURREN(N__27595),
            .RGB2(rgb_b),
            .RGB1PWM(N__19329),
            .RGB0PWM(N__46987),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21300),
            .lcout(pwm_duty_input_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47463),
            .ce(N__24483),
            .sr(N__46905));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_6  (
            .in0(N__19026),
            .in1(N__18293),
            .in2(_gnd_net_),
            .in3(N__18535),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_7_1  (
            .in0(N__18611),
            .in1(N__18266),
            .in2(N__18594),
            .in3(N__18248),
            .lcout(\current_shift_inst.PI_CTRL.m14_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_7_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_7_4  (
            .in0(N__18249),
            .in1(N__18359),
            .in2(N__18452),
            .in3(N__18612),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.m7_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_1_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_1_7_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_1_7_5  (
            .in0(N__18593),
            .in1(N__18536),
            .in2(N__18180),
            .in3(N__18267),
            .lcout(i8_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_0  (
            .in0(N__18325),
            .in1(N__19432),
            .in2(N__20592),
            .in3(N__18313),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47460),
            .ce(N__24465),
            .sr(N__46918));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_8_2 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_8_2  (
            .in0(N__18326),
            .in1(N__19433),
            .in2(N__20898),
            .in3(N__18314),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47460),
            .ce(N__24465),
            .sr(N__46918));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_8_6 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_8_6  (
            .in0(N__18327),
            .in1(N__19434),
            .in2(N__20871),
            .in3(N__18315),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47460),
            .ce(N__24465),
            .sr(N__46918));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__19841),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__18228),
            .in2(_gnd_net_),
            .in3(N__18219),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__18216),
            .in2(_gnd_net_),
            .in3(N__18207),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__18204),
            .in2(_gnd_net_),
            .in3(N__18195),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__18618),
            .in2(_gnd_net_),
            .in3(N__18192),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__27716),
            .in2(N__18936),
            .in3(N__18189),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(N__18894),
            .in2(N__27776),
            .in3(N__18186),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(N__18855),
            .in2(N__27777),
            .in3(N__18183),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__18816),
            .in2(_gnd_net_),
            .in3(N__18231),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__18777),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__18738),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__18699),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__19218),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__19179),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__19152),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__19128),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__19101),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__19077),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__19050),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__18975),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18303),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_11_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_11_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__18671),
            .in2(_gnd_net_),
            .in3(N__19948),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6  (
            .in0(N__18300),
            .in1(N__19025),
            .in2(N__18282),
            .in3(N__18559),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_12_0 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_12_0  (
            .in0(N__19399),
            .in1(N__21293),
            .in2(N__20679),
            .in3(N__20300),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__24500),
            .sr(N__46935));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_1 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_1  (
            .in0(N__19401),
            .in1(N__19301),
            .in2(N__20846),
            .in3(N__19420),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__24500),
            .sr(N__46935));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_12_2 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_12_2  (
            .in0(N__19397),
            .in1(N__21291),
            .in2(N__20763),
            .in3(N__20298),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__24500),
            .sr(N__46935));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_12_4 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_12_4  (
            .in0(N__19398),
            .in1(N__21292),
            .in2(N__20730),
            .in3(N__20299),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__24500),
            .sr(N__46935));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_12_6 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_12_6  (
            .in0(N__19400),
            .in1(N__21294),
            .in2(N__21063),
            .in3(N__20301),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__24500),
            .sr(N__46935));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_13_4 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_13_4  (
            .in0(N__20297),
            .in1(N__19254),
            .in2(N__20811),
            .in3(N__19350),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47439),
            .ce(N__24510),
            .sr(N__46939));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_13_5 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_13_5  (
            .in0(N__19382),
            .in1(N__21295),
            .in2(N__20640),
            .in3(N__20296),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47439),
            .ce(N__24510),
            .sr(N__46939));
    defparam \current_shift_inst.N_22_i_i_LC_1_30_4 .C_ON=1'b0;
    defparam \current_shift_inst.N_22_i_i_LC_1_30_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.N_22_i_i_LC_1_30_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.N_22_i_i_LC_1_30_4  (
            .in0(N__35073),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46986),
            .lcout(N_22_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_7_0 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_7_0  (
            .in0(N__18333),
            .in1(N__18567),
            .in2(N__18555),
            .in3(N__18453),
            .lcout(N_28_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_8_1 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_8_1  (
            .in0(N__18413),
            .in1(N__18395),
            .in2(N__18381),
            .in3(N__18360),
            .lcout(\current_shift_inst.PI_CTRL.N_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_8_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_8_5  (
            .in0(N__21296),
            .in1(N__19395),
            .in2(_gnd_net_),
            .in3(N__19272),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_8_6 .LUT_INIT=16'b0000111100000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_8_6  (
            .in0(N__19396),
            .in1(N__19302),
            .in2(N__20850),
            .in3(N__19431),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_8_7  (
            .in0(N__19811),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19544),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0  (
            .in0(N__20218),
            .in1(N__19526),
            .in2(N__20199),
            .in3(N__19892),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1  (
            .in0(N__20177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18689),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2  (
            .in0(N__18690),
            .in1(N__20163),
            .in2(N__18681),
            .in3(N__19893),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__20077),
            .in2(_gnd_net_),
            .in3(N__19739),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_4  (
            .in0(N__18678),
            .in1(N__19952),
            .in2(N__19926),
            .in3(N__19890),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(N__19775),
            .in2(_gnd_net_),
            .in3(N__18659),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6  (
            .in0(N__18660),
            .in1(N__19761),
            .in2(N__18651),
            .in3(N__19891),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_7  (
            .in0(N__20117),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19508),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__18648),
            .in2(N__18633),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__18966),
            .in2(N__18954),
            .in3(N__18927),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__18924),
            .in2(N__18912),
            .in3(N__18888),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__18885),
            .in2(N__18873),
            .in3(N__18849),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__18846),
            .in2(N__18834),
            .in3(N__18810),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(N__18807),
            .in2(N__18795),
            .in3(N__18771),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(N__18768),
            .in2(N__18756),
            .in3(N__18732),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(N__18729),
            .in2(N__18717),
            .in3(N__18693),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__19248),
            .in2(N__19236),
            .in3(N__19212),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__19209),
            .in2(N__19197),
            .in3(N__19173),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__19013),
            .in2(N__19170),
            .in3(N__19146),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__19143),
            .in2(N__19027),
            .in3(N__19122),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__19017),
            .in2(N__19119),
            .in3(N__19095),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__19092),
            .in2(N__19028),
            .in3(N__19071),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__19021),
            .in2(N__19068),
            .in3(N__19044),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__19041),
            .in2(N__19029),
            .in3(N__18969),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0  (
            .in0(N__19320),
            .in1(N__19314),
            .in2(_gnd_net_),
            .in3(N__19308),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_1  (
            .in0(N__19287),
            .in1(N__20133),
            .in2(N__19305),
            .in3(N__20147),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__20809),
            .in2(_gnd_net_),
            .in3(N__20836),
            .lcout(\current_shift_inst.PI_CTRL.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_4 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_4  (
            .in0(N__21266),
            .in1(N__20810),
            .in2(_gnd_net_),
            .in3(N__19268),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_12_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_12_6  (
            .in0(N__20148),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19286),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__20749),
            .in2(_gnd_net_),
            .in3(N__21059),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_13_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_13_4  (
            .in0(N__20674),
            .in1(N__20722),
            .in2(N__19275),
            .in3(N__20633),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(\current_shift_inst.PI_CTRL.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_13_5 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_13_5  (
            .in0(N__21265),
            .in1(N__20805),
            .in2(N__19257),
            .in3(N__19376),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_13_7 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_13_7  (
            .in0(N__19440),
            .in1(N__19349),
            .in2(N__21284),
            .in3(N__20275),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOLF4_14_LC_2_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOLF4_14_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOLF4_14_LC_2_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOLF4_14_LC_2_14_2  (
            .in0(N__20964),
            .in1(N__21354),
            .in2(N__21330),
            .in3(N__21387),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_14_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_14_3  (
            .in0(N__20031),
            .in1(N__19335),
            .in2(N__19404),
            .in3(N__20232),
            .lcout(\current_shift_inst.PI_CTRL.N_178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_2_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_2_14_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__20626),
            .in2(_gnd_net_),
            .in3(N__21055),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_14_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_14_6  (
            .in0(N__20675),
            .in1(N__20723),
            .in2(N__19353),
            .in3(N__20756),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_15_LC_2_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_15_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_15_LC_2_15_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_15_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__20946),
            .in2(_gnd_net_),
            .in3(N__21144),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_10_LC_2_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_10_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_10_LC_2_15_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_10_LC_2_15_7  (
            .in0(N__21126),
            .in1(N__20334),
            .in2(N__19338),
            .in3(N__21030),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_2_29_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_29_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_29_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_29_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un7_start_stop_0_a3_LC_2_30_7 .C_ON=1'b0;
    defparam \current_shift_inst.un7_start_stop_0_a3_LC_2_30_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un7_start_stop_0_a3_LC_2_30_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \current_shift_inst.un7_start_stop_0_a3_LC_2_30_7  (
            .in0(_gnd_net_),
            .in1(N__35072),
            .in2(_gnd_net_),
            .in3(N__46985),
            .lcout(un7_start_stop_0_a3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_7_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_7_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_7_0 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_3_7_0  (
            .in0(N__20435),
            .in1(N__20550),
            .in2(N__20499),
            .in3(N__19587),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47458),
            .ce(),
            .sr(N__46892));
    defparam \pwm_generator_inst.threshold_0_LC_3_7_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_3_7_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_3_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_3_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19491),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47458),
            .ce(),
            .sr(N__46892));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_7_2 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_7_2 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_3_7_2  (
            .in0(N__20436),
            .in1(N__20551),
            .in2(N__20500),
            .in3(N__19578),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47458),
            .ce(),
            .sr(N__46892));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_7_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_7_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_7_4 .LUT_INIT=16'b0100010000001100;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_3_7_4  (
            .in0(N__20434),
            .in1(N__19479),
            .in2(N__20498),
            .in3(N__20549),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47458),
            .ce(),
            .sr(N__46892));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_7_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_7_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_7_7 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_3_7_7  (
            .in0(N__20548),
            .in1(N__20482),
            .in2(N__20447),
            .in3(N__19449),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47458),
            .ce(),
            .sr(N__46892));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0  (
            .in0(_gnd_net_),
            .in1(N__19485),
            .in2(N__19911),
            .in3(N__19909),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_3_8_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1  (
            .in0(_gnd_net_),
            .in1(N__19827),
            .in2(_gnd_net_),
            .in3(N__19473),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2  (
            .in0(_gnd_net_),
            .in1(N__19533),
            .in2(_gnd_net_),
            .in3(N__19470),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19467),
            .in3(N__19458),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4  (
            .in0(_gnd_net_),
            .in1(N__19455),
            .in2(_gnd_net_),
            .in3(N__19443),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5  (
            .in0(_gnd_net_),
            .in1(N__19608),
            .in2(_gnd_net_),
            .in3(N__19602),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6  (
            .in0(_gnd_net_),
            .in1(N__19599),
            .in2(_gnd_net_),
            .in3(N__19581),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7  (
            .in0(_gnd_net_),
            .in1(N__19497),
            .in2(_gnd_net_),
            .in3(N__19572),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19728),
            .in3(N__19569),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1  (
            .in0(N__19904),
            .in1(N__20040),
            .in2(N__19566),
            .in3(N__19551),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_9_3 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_9_3  (
            .in0(N__19900),
            .in1(N__19548),
            .in2(N__19791),
            .in3(N__19810),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_9_4  (
            .in0(N__20219),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19527),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_9_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_9_7  (
            .in0(N__20097),
            .in1(N__20116),
            .in2(N__19910),
            .in3(N__19512),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_10_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_10_0 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_10_0  (
            .in0(N__19905),
            .in1(N__19746),
            .in2(N__20081),
            .in3(N__20055),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_3_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_3_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_3_10_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_3_10_5  (
            .in0(N__37410),
            .in1(N__40893),
            .in2(_gnd_net_),
            .in3(N__37680),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47447),
            .ce(N__30888),
            .sr(N__46919));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_11_0  (
            .in0(_gnd_net_),
            .in1(N__19707),
            .in2(_gnd_net_),
            .in3(N__19719),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_3_11_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(N__19689),
            .in2(_gnd_net_),
            .in3(N__19701),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__19671),
            .in2(_gnd_net_),
            .in3(N__19683),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(N__19653),
            .in2(_gnd_net_),
            .in3(N__19665),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(N__19632),
            .in2(_gnd_net_),
            .in3(N__19647),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_11_5  (
            .in0(_gnd_net_),
            .in1(N__19614),
            .in2(_gnd_net_),
            .in3(N__19626),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_11_6  (
            .in0(_gnd_net_),
            .in1(N__20013),
            .in2(_gnd_net_),
            .in3(N__20025),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_11_7  (
            .in0(_gnd_net_),
            .in1(N__19995),
            .in2(_gnd_net_),
            .in3(N__20007),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__19977),
            .in2(_gnd_net_),
            .in3(N__19989),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_3_12_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_12_1  (
            .in0(_gnd_net_),
            .in1(N__19959),
            .in2(_gnd_net_),
            .in3(N__19971),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(N__19953),
            .in2(_gnd_net_),
            .in3(N__19914),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_12_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_12_3  (
            .in0(N__19865),
            .in1(N__19845),
            .in2(_gnd_net_),
            .in3(N__19818),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_12_4  (
            .in0(_gnd_net_),
            .in1(N__19815),
            .in2(_gnd_net_),
            .in3(N__19779),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_12_5  (
            .in0(_gnd_net_),
            .in1(N__19776),
            .in2(_gnd_net_),
            .in3(N__19749),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_12_6  (
            .in0(_gnd_net_),
            .in1(N__20220),
            .in2(_gnd_net_),
            .in3(N__20184),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_12_7  (
            .in0(_gnd_net_),
            .in1(N__20181),
            .in2(_gnd_net_),
            .in3(N__20151),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(N__20146),
            .in2(_gnd_net_),
            .in3(N__20127),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_3_13_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20124),
            .in3(N__20085),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(N__20082),
            .in2(_gnd_net_),
            .in3(N__20046),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_13_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20043),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIC5B4_11_LC_3_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIC5B4_11_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIC5B4_11_LC_3_14_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIC5B4_11_LC_3_14_1  (
            .in0(N__20994),
            .in1(N__20925),
            .in2(N__21009),
            .in3(N__20981),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIG72_10_LC_3_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIG72_10_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIG72_10_LC_3_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIG72_10_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__21323),
            .in2(_gnd_net_),
            .in3(N__21023),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRKT8_11_LC_3_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRKT8_11_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRKT8_11_LC_3_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRKT8_11_LC_3_14_4  (
            .in0(N__21386),
            .in1(N__21005),
            .in2(N__20307),
            .in3(N__20247),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_14_5  (
            .in0(N__20241),
            .in1(N__20253),
            .in2(N__20304),
            .in3(N__20259),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3DG5_12_LC_3_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3DG5_12_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3DG5_12_LC_3_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3DG5_12_LC_3_14_7  (
            .in0(N__20993),
            .in1(N__20960),
            .in2(N__21105),
            .in3(N__20226),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_3_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_3_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_3_15_0  (
            .in0(N__21194),
            .in1(N__21206),
            .in2(N__21125),
            .in3(N__20939),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_20_LC_3_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_20_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_20_LC_3_15_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_20_LC_3_15_2  (
            .in0(N__21140),
            .in1(N__21155),
            .in2(N__21350),
            .in3(N__21170),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOJD4_13_LC_3_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOJD4_13_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOJD4_13_LC_3_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOJD4_13_LC_3_15_3  (
            .in0(N__21081),
            .in1(N__20924),
            .in2(N__20982),
            .in3(N__21365),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_3_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_3_15_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__21207),
            .in2(_gnd_net_),
            .in3(N__21171),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_19_LC_3_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_19_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_19_LC_3_15_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_19_LC_3_15_5  (
            .in0(N__21183),
            .in1(N__21366),
            .in2(N__20235),
            .in3(N__21080),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0U62_19_LC_3_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0U62_19_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0U62_19_LC_3_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0U62_19_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__21398),
            .in2(_gnd_net_),
            .in3(N__21182),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_18_LC_3_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_18_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_18_LC_3_15_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_18_LC_3_15_7  (
            .in0(N__21399),
            .in1(N__21101),
            .in2(N__21159),
            .in3(N__21195),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_counter_cry_1_c_LC_4_5_0.C_ON=1'b1;
    defparam un5_counter_cry_1_c_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam un5_counter_cry_1_c_LC_4_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_counter_cry_1_c_LC_4_5_0 (
            .in0(_gnd_net_),
            .in1(N__21581),
            .in2(N__22077),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(un5_counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_2_LC_4_5_1.C_ON=1'b1;
    defparam counter_2_LC_4_5_1.SEQ_MODE=4'b1010;
    defparam counter_2_LC_4_5_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_2_LC_4_5_1 (
            .in0(_gnd_net_),
            .in1(N__21594),
            .in2(_gnd_net_),
            .in3(N__20328),
            .lcout(counterZ0Z_2),
            .ltout(),
            .carryin(un5_counter_cry_1),
            .carryout(un5_counter_cry_2),
            .clk(N__47461),
            .ce(),
            .sr(N__46866));
    defparam counter_3_LC_4_5_2.C_ON=1'b1;
    defparam counter_3_LC_4_5_2.SEQ_MODE=4'b1010;
    defparam counter_3_LC_4_5_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_3_LC_4_5_2 (
            .in0(_gnd_net_),
            .in1(N__21486),
            .in2(_gnd_net_),
            .in3(N__20325),
            .lcout(counterZ0Z_3),
            .ltout(),
            .carryin(un5_counter_cry_2),
            .carryout(un5_counter_cry_3),
            .clk(N__47461),
            .ce(),
            .sr(N__46866));
    defparam counter_4_LC_4_5_3.C_ON=1'b1;
    defparam counter_4_LC_4_5_3.SEQ_MODE=4'b1010;
    defparam counter_4_LC_4_5_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_4_LC_4_5_3 (
            .in0(_gnd_net_),
            .in1(N__21513),
            .in2(_gnd_net_),
            .in3(N__20322),
            .lcout(counterZ0Z_4),
            .ltout(),
            .carryin(un5_counter_cry_3),
            .carryout(un5_counter_cry_4),
            .clk(N__47461),
            .ce(),
            .sr(N__46866));
    defparam counter_5_LC_4_5_4.C_ON=1'b1;
    defparam counter_5_LC_4_5_4.SEQ_MODE=4'b1010;
    defparam counter_5_LC_4_5_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_5_LC_4_5_4 (
            .in0(_gnd_net_),
            .in1(N__21525),
            .in2(_gnd_net_),
            .in3(N__20319),
            .lcout(counterZ0Z_5),
            .ltout(),
            .carryin(un5_counter_cry_4),
            .carryout(un5_counter_cry_5),
            .clk(N__47461),
            .ce(),
            .sr(N__46866));
    defparam counter_6_LC_4_5_5.C_ON=1'b1;
    defparam counter_6_LC_4_5_5.SEQ_MODE=4'b1010;
    defparam counter_6_LC_4_5_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_6_LC_4_5_5 (
            .in0(_gnd_net_),
            .in1(N__21500),
            .in2(_gnd_net_),
            .in3(N__20316),
            .lcout(counterZ0Z_6),
            .ltout(),
            .carryin(un5_counter_cry_5),
            .carryout(un5_counter_cry_6),
            .clk(N__47461),
            .ce(),
            .sr(N__46866));
    defparam counter_RNO_0_7_LC_4_5_6.C_ON=1'b1;
    defparam counter_RNO_0_7_LC_4_5_6.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_7_LC_4_5_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_7_LC_4_5_6 (
            .in0(_gnd_net_),
            .in1(N__21219),
            .in2(_gnd_net_),
            .in3(N__20313),
            .lcout(counter_RNO_0Z0Z_7),
            .ltout(),
            .carryin(un5_counter_cry_6),
            .carryout(un5_counter_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_8_LC_4_5_7.C_ON=1'b1;
    defparam counter_8_LC_4_5_7.SEQ_MODE=4'b1010;
    defparam counter_8_LC_4_5_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_8_LC_4_5_7 (
            .in0(_gnd_net_),
            .in1(N__21561),
            .in2(_gnd_net_),
            .in3(N__20310),
            .lcout(counterZ0Z_8),
            .ltout(),
            .carryin(un5_counter_cry_7),
            .carryout(un5_counter_cry_8),
            .clk(N__47461),
            .ce(),
            .sr(N__46866));
    defparam counter_9_LC_4_6_0.C_ON=1'b1;
    defparam counter_9_LC_4_6_0.SEQ_MODE=4'b1010;
    defparam counter_9_LC_4_6_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_9_LC_4_6_0 (
            .in0(_gnd_net_),
            .in1(N__21537),
            .in2(_gnd_net_),
            .in3(N__20370),
            .lcout(counterZ0Z_9),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(un5_counter_cry_9),
            .clk(N__47459),
            .ce(),
            .sr(N__46876));
    defparam counter_RNO_0_10_LC_4_6_1.C_ON=1'b1;
    defparam counter_RNO_0_10_LC_4_6_1.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_10_LC_4_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_10_LC_4_6_1 (
            .in0(_gnd_net_),
            .in1(N__21411),
            .in2(_gnd_net_),
            .in3(N__20367),
            .lcout(counter_RNO_0Z0Z_10),
            .ltout(),
            .carryin(un5_counter_cry_9),
            .carryout(un5_counter_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_11_LC_4_6_2.C_ON=1'b1;
    defparam counter_11_LC_4_6_2.SEQ_MODE=4'b1010;
    defparam counter_11_LC_4_6_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_11_LC_4_6_2 (
            .in0(_gnd_net_),
            .in1(N__21549),
            .in2(_gnd_net_),
            .in3(N__20364),
            .lcout(counterZ0Z_11),
            .ltout(),
            .carryin(un5_counter_cry_10),
            .carryout(un5_counter_cry_11),
            .clk(N__47459),
            .ce(),
            .sr(N__46876));
    defparam counter_RNO_0_12_LC_4_6_3.C_ON=1'b0;
    defparam counter_RNO_0_12_LC_4_6_3.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_12_LC_4_6_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 counter_RNO_0_12_LC_4_6_3 (
            .in0(_gnd_net_),
            .in1(N__21434),
            .in2(_gnd_net_),
            .in3(N__20361),
            .lcout(counter_RNO_0Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_4_7_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_4_7_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_4_7_1 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_4_7_1  (
            .in0(N__20552),
            .in1(N__20490),
            .in2(N__20444),
            .in3(N__20358),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47453),
            .ce(),
            .sr(N__46885));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_7_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_7_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_7_3 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_4_7_3  (
            .in0(N__20553),
            .in1(N__20491),
            .in2(N__20445),
            .in3(N__20352),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47453),
            .ce(),
            .sr(N__46885));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_7_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_7_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_7_4 .LUT_INIT=16'b1111111111001010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_4_7_4  (
            .in0(N__20489),
            .in1(N__20424),
            .in2(N__20563),
            .in3(N__20346),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47453),
            .ce(),
            .sr(N__46885));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_7_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_7_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_7_7 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_4_7_7  (
            .in0(N__20554),
            .in1(N__20492),
            .in2(N__20446),
            .in3(N__20340),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47453),
            .ce(),
            .sr(N__46885));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25344),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47451),
            .ce(N__24466),
            .sr(N__46893));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_4_8_7  (
            .in0(N__25284),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47451),
            .ce(N__24466),
            .sr(N__46893));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_9_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_9_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_9_0 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_4_9_0  (
            .in0(N__20501),
            .in1(N__20565),
            .in2(N__20574),
            .in3(N__20440),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__46906));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_4_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_4_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_4_9_1 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_4_9_1  (
            .in0(N__20564),
            .in1(N__20502),
            .in2(N__20448),
            .in3(N__20382),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__46906));
    defparam \pwm_generator_inst.threshold_9_LC_4_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_4_9_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_4_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20376),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__46906));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_4_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_4_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_4_10_0 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_4_10_0  (
            .in0(N__24653),
            .in1(N__21672),
            .in2(N__24885),
            .in3(N__24977),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__24485),
            .sr(N__46912));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_4_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_4_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_4_10_1 .LUT_INIT=16'b1100110100001101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_4_10_1  (
            .in0(N__24978),
            .in1(N__21663),
            .in2(N__24890),
            .in3(N__24654),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__24485),
            .sr(N__46912));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_10_2 .LUT_INIT=16'b1000110010001111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_4_10_2  (
            .in0(N__24655),
            .in1(N__21654),
            .in2(N__24886),
            .in3(N__24979),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__24485),
            .sr(N__46912));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_4_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_4_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_4_10_3 .LUT_INIT=16'b1100110100001101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_4_10_3  (
            .in0(N__24980),
            .in1(N__21645),
            .in2(N__24891),
            .in3(N__24656),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__24485),
            .sr(N__46912));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_10_4 .LUT_INIT=16'b1000110010001111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_4_10_4  (
            .in0(N__24657),
            .in1(N__21834),
            .in2(N__24887),
            .in3(N__24981),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__24485),
            .sr(N__46912));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_4_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_4_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_4_10_5 .LUT_INIT=16'b1111000100110001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_4_10_5  (
            .in0(N__24982),
            .in1(N__24840),
            .in2(N__21825),
            .in3(N__24658),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__24485),
            .sr(N__46912));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_4_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_4_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_4_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24257),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__24485),
            .sr(N__46912));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_4_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_4_11_0 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_4_11_0  (
            .in0(N__21698),
            .in1(N__21721),
            .in2(N__22528),
            .in3(N__21745),
            .lcout(\current_shift_inst.PI_CTRL.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_4_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_4_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_4_11_5 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_4_11_5  (
            .in0(N__21942),
            .in1(N__24659),
            .in2(N__24892),
            .in3(N__25023),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47431),
            .ce(N__24492),
            .sr(N__46920));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_4_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_4_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_4_12_0 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_4_12_0  (
            .in0(N__24662),
            .in1(N__21861),
            .in2(N__24889),
            .in3(N__25026),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47424),
            .ce(N__24468),
            .sr(N__46924));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24282),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47424),
            .ce(N__24468),
            .sr(N__46924));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_4_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_4_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_4_12_2 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_4_12_2  (
            .in0(N__24660),
            .in1(N__21882),
            .in2(N__24888),
            .in3(N__25024),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47424),
            .ce(N__24468),
            .sr(N__46924));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_4_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_4_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_4_12_3 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_4_12_3  (
            .in0(N__25025),
            .in1(N__24850),
            .in2(N__21873),
            .in3(N__24661),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47424),
            .ce(N__24468),
            .sr(N__46924));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_4_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_4_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_4_12_5 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_4_12_5  (
            .in0(N__25027),
            .in1(N__24851),
            .in2(N__21852),
            .in3(N__24663),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47424),
            .ce(N__24468),
            .sr(N__46924));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_4_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_4_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_4_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24234),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47424),
            .ce(N__24468),
            .sr(N__46924));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__21753),
            .in2(N__20604),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__47416),
            .ce(N__24502),
            .sr(N__46927));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__21729),
            .in2(N__20910),
            .in3(N__20880),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__47416),
            .ce(N__24502),
            .sr(N__46927));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__20877),
            .in2(N__21702),
            .in3(N__20853),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__47416),
            .ce(N__24502),
            .sr(N__46927));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__22533),
            .in2(N__22152),
            .in3(N__20814),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__47416),
            .ce(N__24502),
            .sr(N__46927));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__22566),
            .in2(N__22881),
            .in3(N__20775),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__47416),
            .ce(N__24502),
            .sr(N__46927));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(N__20772),
            .in2(N__22374),
            .in3(N__20733),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__47416),
            .ce(N__24502),
            .sr(N__46927));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__22404),
            .in2(N__21909),
            .in3(N__20697),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__47416),
            .ce(N__24502),
            .sr(N__46927));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__22433),
            .in2(N__20694),
            .in3(N__20643),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__47416),
            .ce(N__24502),
            .sr(N__46927));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__22491),
            .in2(N__22128),
            .in3(N__20607),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__47408),
            .ce(N__24507),
            .sr(N__46931));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__21606),
            .in2(N__22464),
            .in3(N__21033),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__47408),
            .ce(N__24507),
            .sr(N__46931));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__22038),
            .in2(N__25077),
            .in3(N__21012),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__47408),
            .ce(N__24507),
            .sr(N__46931));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__23145),
            .in2(N__22113),
            .in3(N__20997),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__47408),
            .ce(N__24507),
            .sr(N__46931));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__22697),
            .in2(N__22023),
            .in3(N__20985),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__47408),
            .ce(N__24507),
            .sr(N__46931));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(N__23226),
            .in2(N__22032),
            .in3(N__20967),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__47408),
            .ce(N__24507),
            .sr(N__46931));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(N__23250),
            .in2(N__21921),
            .in3(N__20949),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__47408),
            .ce(N__24507),
            .sr(N__46931));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(N__22617),
            .in2(N__22008),
            .in3(N__20928),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__47408),
            .ce(N__24507),
            .sr(N__46931));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__21999),
            .in2(N__23190),
            .in3(N__20913),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__47399),
            .ce(N__24508),
            .sr(N__46936));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__24540),
            .in2(N__21981),
            .in3(N__21198),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__47399),
            .ce(N__24508),
            .sr(N__46936));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__23964),
            .in2(N__21993),
            .in3(N__21186),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__47399),
            .ce(N__24508),
            .sr(N__46936));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__23106),
            .in2(N__22137),
            .in3(N__21174),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__47399),
            .ce(N__24508),
            .sr(N__46936));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__23074),
            .in2(N__21960),
            .in3(N__21162),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__47399),
            .ce(N__24508),
            .sr(N__46936));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__23822),
            .in2(N__25110),
            .in3(N__21147),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__47399),
            .ce(N__24508),
            .sr(N__46936));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(N__23045),
            .in2(N__22101),
            .in3(N__21129),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__47399),
            .ce(N__24508),
            .sr(N__46936));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__22083),
            .in2(N__22647),
            .in3(N__21108),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__47399),
            .ce(N__24508),
            .sr(N__46936));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__23859),
            .in2(N__22092),
            .in3(N__21084),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__47389),
            .ce(N__24509),
            .sr(N__46940));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__22917),
            .in2(N__23904),
            .in3(N__21066),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__47389),
            .ce(N__24509),
            .sr(N__46940));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__22925),
            .in2(N__23787),
            .in3(N__21390),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__47389),
            .ce(N__24509),
            .sr(N__46940));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__22856),
            .in2(N__22934),
            .in3(N__21369),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__47389),
            .ce(N__24509),
            .sr(N__46940));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__22736),
            .in2(N__22932),
            .in3(N__21357),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__47389),
            .ce(N__24509),
            .sr(N__46940));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(N__23292),
            .in2(N__22935),
            .in3(N__21333),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__47389),
            .ce(N__24509),
            .sr(N__46940));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__22983),
            .in2(N__22933),
            .in3(N__21306),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__47389),
            .ce(N__24509),
            .sr(N__46940));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7  (
            .in0(N__24867),
            .in1(N__22924),
            .in2(_gnd_net_),
            .in3(N__21303),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47389),
            .ce(N__24509),
            .sr(N__46940));
    defparam counter_7_LC_5_4_0.C_ON=1'b0;
    defparam counter_7_LC_5_4_0.SEQ_MODE=4'b1010;
    defparam counter_7_LC_5_4_0.LUT_INIT=16'b0111000011110000;
    LogicCell40 counter_7_LC_5_4_0 (
            .in0(N__22314),
            .in1(N__22272),
            .in2(N__21228),
            .in3(N__22227),
            .lcout(counterZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47462),
            .ce(),
            .sr(N__46848));
    defparam counter_1_LC_5_4_1.C_ON=1'b0;
    defparam counter_1_LC_5_4_1.SEQ_MODE=4'b1010;
    defparam counter_1_LC_5_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_1_LC_5_4_1 (
            .in0(_gnd_net_),
            .in1(N__21582),
            .in2(_gnd_net_),
            .in3(N__22072),
            .lcout(counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47462),
            .ce(),
            .sr(N__46848));
    defparam counter_RNI800G_7_LC_5_5_2.C_ON=1'b0;
    defparam counter_RNI800G_7_LC_5_5_2.SEQ_MODE=4'b0000;
    defparam counter_RNI800G_7_LC_5_5_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 counter_RNI800G_7_LC_5_5_2 (
            .in0(_gnd_net_),
            .in1(N__21410),
            .in2(_gnd_net_),
            .in3(N__21218),
            .lcout(),
            .ltout(un2_counter_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI3BSP_1_LC_5_5_3.C_ON=1'b0;
    defparam counter_RNI3BSP_1_LC_5_5_3.SEQ_MODE=4'b0000;
    defparam counter_RNI3BSP_1_LC_5_5_3.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNI3BSP_1_LC_5_5_3 (
            .in0(N__21593),
            .in1(N__21580),
            .in2(N__21564),
            .in3(N__22073),
            .lcout(un2_counter_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIM6001_12_LC_5_5_4.C_ON=1'b0;
    defparam counter_RNIM6001_12_LC_5_5_4.SEQ_MODE=4'b0000;
    defparam counter_RNIM6001_12_LC_5_5_4.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNIM6001_12_LC_5_5_4 (
            .in0(N__21560),
            .in1(N__21548),
            .in2(N__21435),
            .in3(N__21536),
            .lcout(un2_counter_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNII76D_3_LC_5_5_5.C_ON=1'b0;
    defparam counter_RNII76D_3_LC_5_5_5.SEQ_MODE=4'b0000;
    defparam counter_RNII76D_3_LC_5_5_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 counter_RNII76D_3_LC_5_5_5 (
            .in0(N__21524),
            .in1(N__21512),
            .in2(N__21501),
            .in3(N__21485),
            .lcout(un2_counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_4_LC_5_6_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_5_6_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_5_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21474),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(),
            .sr(N__46867));
    defparam \pwm_generator_inst.threshold_2_LC_5_6_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_5_6_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_5_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21462),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(),
            .sr(N__46867));
    defparam \pwm_generator_inst.threshold_6_LC_5_6_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_5_6_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_5_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21456),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(),
            .sr(N__46867));
    defparam counter_12_LC_5_6_5.C_ON=1'b0;
    defparam counter_12_LC_5_6_5.SEQ_MODE=4'b1010;
    defparam counter_12_LC_5_6_5.LUT_INIT=16'b0111000011110000;
    LogicCell40 counter_12_LC_5_6_5 (
            .in0(N__22313),
            .in1(N__22271),
            .in2(N__21444),
            .in3(N__22226),
            .lcout(counterZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(),
            .sr(N__46867));
    defparam counter_10_LC_5_6_7.C_ON=1'b0;
    defparam counter_10_LC_5_6_7.SEQ_MODE=4'b1010;
    defparam counter_10_LC_5_6_7.LUT_INIT=16'b0111000011110000;
    LogicCell40 counter_10_LC_5_6_7 (
            .in0(N__22312),
            .in1(N__22270),
            .in2(N__21420),
            .in3(N__22225),
            .lcout(counterZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(),
            .sr(N__46867));
    defparam \pwm_generator_inst.threshold_8_LC_5_7_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_5_7_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_5_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21636),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47452),
            .ce(),
            .sr(N__46877));
    defparam \pwm_generator_inst.threshold_3_LC_5_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_5_7_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_5_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21627),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47452),
            .ce(),
            .sr(N__46877));
    defparam \pwm_generator_inst.threshold_7_LC_5_7_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_5_7_3 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_5_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21621),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47452),
            .ce(),
            .sr(N__46877));
    defparam \pwm_generator_inst.threshold_5_LC_5_7_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_5_7_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_5_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_5_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21612),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47452),
            .ce(),
            .sr(N__46877));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25224),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47449),
            .ce(N__24407),
            .sr(N__46886));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_5_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_5_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_5_9_0 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_5_9_0  (
            .in0(N__24605),
            .in1(N__21894),
            .in2(N__24897),
            .in3(N__25005),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47441),
            .ce(N__24475),
            .sr(N__46894));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_5_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_5_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_5_9_2 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_5_9_2  (
            .in0(N__24604),
            .in1(N__21765),
            .in2(N__24896),
            .in3(N__25004),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47441),
            .ce(N__24475),
            .sr(N__46894));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4  (
            .in0(N__24601),
            .in1(N__21810),
            .in2(N__24894),
            .in3(N__25001),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47441),
            .ce(N__24475),
            .sr(N__46894));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_5_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_5_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_5_9_6 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_5_9_6  (
            .in0(N__24602),
            .in1(N__21798),
            .in2(N__24895),
            .in3(N__25002),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47441),
            .ce(N__24475),
            .sr(N__46894));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_5_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_5_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_5_9_7 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_5_9_7  (
            .in0(N__25003),
            .in1(N__24872),
            .in2(N__21786),
            .in3(N__24603),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47441),
            .ce(N__24475),
            .sr(N__46894));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_5_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_5_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_5_10_0 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__21746),
            .in2(N__24281),
            .in3(N__22802),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .clk(N__47432),
            .ce(N__24484),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_5_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_5_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_5_10_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_5_10_1  (
            .in0(N__22800),
            .in1(N__21722),
            .in2(N__24258),
            .in3(N__21705),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(N__47432),
            .ce(N__24484),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_5_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_5_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_5_10_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_5_10_2  (
            .in0(N__22803),
            .in1(N__21697),
            .in2(N__24233),
            .in3(N__21678),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(N__47432),
            .ce(N__24484),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_5_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_5_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_5_10_3 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_5_10_3  (
            .in0(N__22801),
            .in1(N__22527),
            .in2(N__24207),
            .in3(N__21675),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(N__47432),
            .ce(N__24484),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_5_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_5_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__22560),
            .in2(N__25368),
            .in3(N__21666),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_5_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_5_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(N__22357),
            .in2(N__25343),
            .in3(N__21657),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_5_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_5_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(N__22398),
            .in2(N__25311),
            .in3(N__21648),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_5_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_5_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__22425),
            .in2(N__25283),
            .in3(N__21639),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_5_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_5_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__22485),
            .in2(N__25254),
            .in3(N__21828),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_5_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__22455),
            .in2(N__25223),
            .in3(N__21816),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_5_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__25191),
            .in2(N__25076),
            .in3(N__21813),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_5_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__25166),
            .in2(N__23144),
            .in3(N__21801),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_5_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__25595),
            .in2(N__22696),
            .in3(N__21789),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_5_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_5_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__23220),
            .in2(N__25575),
            .in3(N__21774),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_5_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_5_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__23257),
            .in2(N__25551),
            .in3(N__21771),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_5_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_5_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__22613),
            .in2(N__25527),
            .in3(N__21768),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_5_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_5_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__23175),
            .in2(N__25503),
            .in3(N__21756),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_5_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_5_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__24536),
            .in2(N__25476),
            .in3(N__21897),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_5_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_5_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__23944),
            .in2(N__25449),
            .in3(N__21885),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_5_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_5_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__23100),
            .in2(N__25419),
            .in3(N__21876),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_5_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_5_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__23073),
            .in2(N__25392),
            .in3(N__21864),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_5_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_5_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__23808),
            .in2(N__25737),
            .in3(N__21855),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_5_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_5_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__23037),
            .in2(N__25710),
            .in3(N__21843),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_5_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_5_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__22643),
            .in2(N__25683),
            .in3(N__21840),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_5_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_5_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__23855),
            .in2(N__25656),
            .in3(N__21837),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_5_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_5_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__27221),
            .in2(N__23898),
            .in3(N__21951),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_5_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_5_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__23779),
            .in2(N__27237),
            .in3(N__21948),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_5_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_5_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__27225),
            .in2(N__22857),
            .in3(N__21945),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_5_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_5_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__22735),
            .in2(N__27238),
            .in3(N__21933),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_5_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_5_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__23288),
            .in2(N__27243),
            .in3(N__21930),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_5_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_5_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__22978),
            .in2(N__27239),
            .in3(N__21927),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_5_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_5_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_5_13_7  (
            .in0(N__24782),
            .in1(N__27232),
            .in2(_gnd_net_),
            .in3(N__21924),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25550),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47400),
            .ce(N__24506),
            .sr(N__46928));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25310),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47400),
            .ce(N__24506),
            .sr(N__46928));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25190),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47400),
            .ce(N__24506),
            .sr(N__46928));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25574),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47400),
            .ce(N__24506),
            .sr(N__46928));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25596),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47400),
            .ce(N__24506),
            .sr(N__46928));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_5_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_5_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_5_14_5 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_5_14_5  (
            .in0(N__22014),
            .in1(N__24671),
            .in2(N__24871),
            .in3(N__25034),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47400),
            .ce(N__24506),
            .sr(N__46928));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_7  (
            .in0(N__25526),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47400),
            .ce(N__24506),
            .sr(N__46928));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25499),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47390),
            .ce(N__24499),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25442),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47390),
            .ce(N__24499),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25472),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47390),
            .ce(N__24499),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_5_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_5_15_4 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_5_15_4  (
            .in0(N__21969),
            .in1(N__24672),
            .in2(N__24893),
            .in3(N__25035),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47390),
            .ce(N__24499),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_5_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_5_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_5_15_5  (
            .in0(N__25388),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47390),
            .ce(N__24499),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24206),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47390),
            .ce(N__24499),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25415),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47390),
            .ce(N__24499),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25253),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47381),
            .ce(N__24501),
            .sr(N__46937));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25167),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47381),
            .ce(N__24501),
            .sr(N__46937));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25709),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47381),
            .ce(N__24501),
            .sr(N__46937));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25652),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47381),
            .ce(N__24501),
            .sr(N__46937));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25682),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47381),
            .ce(N__24501),
            .sr(N__46937));
    defparam counter_0_LC_7_4_1.C_ON=1'b0;
    defparam counter_0_LC_7_4_1.SEQ_MODE=4'b1010;
    defparam counter_0_LC_7_4_1.LUT_INIT=16'b0000011100001111;
    LogicCell40 counter_0_LC_7_4_1 (
            .in0(N__22236),
            .in1(N__22329),
            .in2(N__22071),
            .in3(N__22283),
            .lcout(counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47455),
            .ce(),
            .sr(N__46836));
    defparam clk_10khz_RNIIENA2_LC_7_5_2.C_ON=1'b0;
    defparam clk_10khz_RNIIENA2_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam clk_10khz_RNIIENA2_LC_7_5_2.LUT_INIT=16'b0111100011110000;
    LogicCell40 clk_10khz_RNIIENA2_LC_7_5_2 (
            .in0(N__22321),
            .in1(N__22273),
            .in2(N__22194),
            .in3(N__22228),
            .lcout(clk_10khz_RNIIENAZ0Z2),
            .ltout(clk_10khz_RNIIENAZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_7_5_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_7_5_3 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_7_5_3  (
            .in0(N__35047),
            .in1(_gnd_net_),
            .in2(N__22338),
            .in3(N__22191),
            .lcout(N_655_g),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_7_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_7_6_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \current_shift_inst.phase_valid_RNISLOR2_LC_7_6_5  (
            .in0(N__28998),
            .in1(N__22192),
            .in2(N__35059),
            .in3(N__22335),
            .lcout(\current_shift_inst.phase_valid_RNISLORZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_10khz_LC_7_6_7.C_ON=1'b0;
    defparam clk_10khz_LC_7_6_7.SEQ_MODE=4'b1010;
    defparam clk_10khz_LC_7_6_7.LUT_INIT=16'b0110110011001100;
    LogicCell40 clk_10khz_LC_7_6_7 (
            .in0(N__22328),
            .in1(N__22193),
            .in2(N__22284),
            .in3(N__22235),
            .lcout(clk_10khz_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47450),
            .ce(),
            .sr(N__46849));
    defparam \pwm_generator_inst.threshold_1_LC_7_7_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_7_7_3 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_7_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22173),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47442),
            .ce(),
            .sr(N__46857));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_7_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_7_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__23605),
            .in2(_gnd_net_),
            .in3(N__23653),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_7_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_7_8_2 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_7_8_2  (
            .in0(N__24178),
            .in1(N__23584),
            .in2(N__22164),
            .in3(N__23632),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_7_8_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_7_8_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_7_8_3  (
            .in0(N__22158),
            .in1(N__24131),
            .in2(N__22161),
            .in3(N__24155),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_7_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_7_8_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_7_8_5  (
            .in0(N__24079),
            .in1(N__24010),
            .in2(_gnd_net_),
            .in3(N__24106),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_9_0  (
            .in0(N__22779),
            .in1(N__22584),
            .in2(N__22770),
            .in3(N__22656),
            .lcout(\current_shift_inst.PI_CTRL.N_46_21 ),
            .ltout(\current_shift_inst.PI_CTRL.N_46_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_9_1  (
            .in0(N__23016),
            .in1(N__23961),
            .in2(N__22587),
            .in3(N__22500),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_9_2  (
            .in0(N__23262),
            .in1(N__23224),
            .in2(N__23188),
            .in3(N__23142),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_4_LC_7_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_4_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_4_LC_7_10_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_4_LC_7_10_0  (
            .in0(N__22565),
            .in1(N__22578),
            .in2(_gnd_net_),
            .in3(N__22344),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_10_1  (
            .in0(N__22457),
            .in1(N__22402),
            .in2(N__22434),
            .in3(N__22367),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_10_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_10_2  (
            .in0(N__22490),
            .in1(N__22564),
            .in2(N__22536),
            .in3(N__22529),
            .lcout(\current_shift_inst.PI_CTRL.N_44 ),
            .ltout(\current_shift_inst.PI_CTRL.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_10_3  (
            .in0(N__24823),
            .in1(N__23951),
            .in2(N__22494),
            .in3(N__23015),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_10_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_10_4  (
            .in0(N__22489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22456),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_10_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_10_5  (
            .in0(N__22432),
            .in1(N__22403),
            .in2(N__22377),
            .in3(N__22366),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_10_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_10_6  (
            .in0(N__23993),
            .in1(N__24824),
            .in2(N__23962),
            .in3(N__25121),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_10_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_10_7  (
            .in0(N__22818),
            .in1(N__22812),
            .in2(N__22806),
            .in3(N__23975),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_11_2  (
            .in0(N__22734),
            .in1(N__22846),
            .in2(N__22982),
            .in3(N__22698),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_11_3  (
            .in0(N__23902),
            .in1(N__23854),
            .in2(N__23783),
            .in3(N__23818),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_7_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_7_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_7_11_4 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_7_11_4  (
            .in0(N__22758),
            .in1(N__24641),
            .in2(N__24828),
            .in3(N__24949),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47409),
            .ce(N__24411),
            .sr(N__46895));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_11_5 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_7_11_5  (
            .in0(N__24950),
            .in1(N__24778),
            .in2(N__24670),
            .in3(N__22749),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47409),
            .ce(N__24411),
            .sr(N__46895));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_12_1  (
            .in0(N__22737),
            .in1(N__22842),
            .in2(N__22974),
            .in3(N__22695),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_12_2  (
            .in0(N__25056),
            .in1(N__23280),
            .in2(N__22612),
            .in3(N__22631),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_7_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_7_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_7_12_3  (
            .in0(N__22630),
            .in1(N__22602),
            .in2(N__23287),
            .in3(N__25057),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_12_4  (
            .in0(N__23258),
            .in1(N__23225),
            .in2(N__23189),
            .in3(N__23143),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_12_6  (
            .in0(N__24535),
            .in1(N__23044),
            .in2(N__23079),
            .in3(N__23105),
            .lcout(\current_shift_inst.PI_CTRL.N_47_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_12_7  (
            .in0(N__23104),
            .in1(N__23075),
            .in2(N__23046),
            .in3(N__24534),
            .lcout(\current_shift_inst.PI_CTRL.N_46_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_7_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_7_13_0 .LUT_INIT=16'b1111010011000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_7_13_0  (
            .in0(N__24649),
            .in1(N__24752),
            .in2(N__22998),
            .in3(N__24975),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(N__24476),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_13_1 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_7_13_1  (
            .in0(N__24972),
            .in1(N__22944),
            .in2(N__24819),
            .in3(N__24646),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(N__24476),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_7_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_7_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27233),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(N__24476),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_7_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_7_13_3 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_7_13_3  (
            .in0(N__24971),
            .in1(N__22890),
            .in2(N__24818),
            .in3(N__24645),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(N__24476),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_7_13_4  (
            .in0(N__25361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(N__24476),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_13_5 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_7_13_5  (
            .in0(N__24973),
            .in1(N__22866),
            .in2(N__24820),
            .in3(N__24647),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(N__24476),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_7_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_7_13_6 .LUT_INIT=16'b1111010011000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_7_13_6  (
            .in0(N__24650),
            .in1(N__24753),
            .in2(N__23316),
            .in3(N__24976),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(N__24476),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_7_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_7_13_7 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_7_13_7  (
            .in0(N__24974),
            .in1(N__23301),
            .in2(N__24821),
            .in3(N__24648),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(N__24476),
            .sr(N__46913));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_7_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_7_14_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_7_14_0  (
            .in0(N__28048),
            .in1(N__28414),
            .in2(N__29529),
            .in3(N__29482),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_7_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_7_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__27304),
            .in2(_gnd_net_),
            .in3(N__29635),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_7_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_7_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__29605),
            .in2(_gnd_net_),
            .in3(N__28262),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNILORI_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_7_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_7_14_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_7_14_3  (
            .in0(N__27336),
            .in1(N__27305),
            .in2(N__29673),
            .in3(N__29636),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_7_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_7_14_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__29668),
            .in2(_gnd_net_),
            .in3(N__27335),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_7_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_7_14_5 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_7_14_5  (
            .in0(N__28261),
            .in1(N__29637),
            .in2(N__29607),
            .in3(N__27306),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_7_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_7_14_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_7_14_7  (
            .in0(N__27334),
            .in1(N__28159),
            .in2(N__29718),
            .in3(N__29672),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_7_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_7_15_0 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_7_15_0  (
            .in0(N__29832),
            .in1(N__27408),
            .in2(N__27381),
            .in3(N__29801),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_7_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_7_15_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_7_15_1  (
            .in0(N__27406),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29831),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_7_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_7_15_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_7_15_2  (
            .in0(N__27379),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29800),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_7_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_7_15_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_7_15_3  (
            .in0(N__27407),
            .in1(N__27437),
            .in2(N__29865),
            .in3(N__29830),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_7_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_7_15_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27438),
            .in3(N__29860),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_7_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_7_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_7_15_5  (
            .in0(N__27380),
            .in1(N__30346),
            .in2(N__29805),
            .in3(N__30289),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_7_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_7_15_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_7_15_6  (
            .in0(N__30290),
            .in1(_gnd_net_),
            .in2(N__30351),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_7_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_7_15_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_7_15_7  (
            .in0(N__29861),
            .in1(N__27471),
            .in2(N__29907),
            .in3(N__27433),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_7_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_7_16_0 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_7_16_0  (
            .in0(N__27466),
            .in1(N__29902),
            .in2(N__29949),
            .in3(N__28345),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_7_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_7_16_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_7_16_1  (
            .in0(N__29903),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27467),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_7_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_7_16_2 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_7_16_2  (
            .in0(N__30402),
            .in1(N__27940),
            .in2(N__30203),
            .in3(N__30441),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27945),
            .in3(N__30196),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_7_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_7_16_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_7_16_4  (
            .in0(N__27913),
            .in1(N__27944),
            .in2(N__30204),
            .in3(N__30166),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5  (
            .in0(N__30167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27914),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_6 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_6  (
            .in0(N__27915),
            .in1(N__30137),
            .in2(N__27888),
            .in3(N__30168),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7  (
            .in0(N__30138),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27887),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_17_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_17_7  (
            .in0(N__26969),
            .in1(N__30524),
            .in2(_gnd_net_),
            .in3(N__30477),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.counter_0_LC_7_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_0_LC_7_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_0_LC_7_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_0_LC_7_19_0  (
            .in0(N__26585),
            .in1(N__28648),
            .in2(_gnd_net_),
            .in3(N__23325),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_0 ),
            .clk(N__47345),
            .ce(N__33641),
            .sr(N__46941));
    defparam \current_shift_inst.timer_phase.counter_1_LC_7_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_1_LC_7_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_1_LC_7_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_1_LC_7_19_1  (
            .in0(N__26580),
            .in1(N__28687),
            .in2(_gnd_net_),
            .in3(N__23322),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_1 ),
            .clk(N__47345),
            .ce(N__33641),
            .sr(N__46941));
    defparam \current_shift_inst.timer_phase.counter_2_LC_7_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_2_LC_7_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_2_LC_7_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_2_LC_7_19_2  (
            .in0(N__26586),
            .in1(N__25615),
            .in2(_gnd_net_),
            .in3(N__23319),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_2 ),
            .clk(N__47345),
            .ce(N__33641),
            .sr(N__46941));
    defparam \current_shift_inst.timer_phase.counter_3_LC_7_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_3_LC_7_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_3_LC_7_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_3_LC_7_19_3  (
            .in0(N__26581),
            .in1(N__25975),
            .in2(_gnd_net_),
            .in3(N__23352),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_3 ),
            .clk(N__47345),
            .ce(N__33641),
            .sr(N__46941));
    defparam \current_shift_inst.timer_phase.counter_4_LC_7_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_4_LC_7_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_4_LC_7_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_4_LC_7_19_4  (
            .in0(N__26587),
            .in1(N__25949),
            .in2(_gnd_net_),
            .in3(N__23349),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_4 ),
            .clk(N__47345),
            .ce(N__33641),
            .sr(N__46941));
    defparam \current_shift_inst.timer_phase.counter_5_LC_7_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_5_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_5_LC_7_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_5_LC_7_19_5  (
            .in0(N__26582),
            .in1(N__25930),
            .in2(_gnd_net_),
            .in3(N__23346),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_5 ),
            .clk(N__47345),
            .ce(N__33641),
            .sr(N__46941));
    defparam \current_shift_inst.timer_phase.counter_6_LC_7_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_6_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_6_LC_7_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_6_LC_7_19_6  (
            .in0(N__26584),
            .in1(N__25898),
            .in2(_gnd_net_),
            .in3(N__23343),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_6 ),
            .clk(N__47345),
            .ce(N__33641),
            .sr(N__46941));
    defparam \current_shift_inst.timer_phase.counter_7_LC_7_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_7_LC_7_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_7_LC_7_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_7_LC_7_19_7  (
            .in0(N__26583),
            .in1(N__25868),
            .in2(_gnd_net_),
            .in3(N__23340),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_7 ),
            .clk(N__47345),
            .ce(N__33641),
            .sr(N__46941));
    defparam \current_shift_inst.timer_phase.counter_8_LC_7_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_8_LC_7_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_8_LC_7_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_8_LC_7_20_0  (
            .in0(N__26591),
            .in1(N__25843),
            .in2(_gnd_net_),
            .in3(N__23337),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_8 ),
            .clk(N__47337),
            .ce(N__33645),
            .sr(N__46943));
    defparam \current_shift_inst.timer_phase.counter_9_LC_7_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_9_LC_7_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_9_LC_7_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_9_LC_7_20_1  (
            .in0(N__26595),
            .in1(N__25813),
            .in2(_gnd_net_),
            .in3(N__23334),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_9 ),
            .clk(N__47337),
            .ce(N__33645),
            .sr(N__46943));
    defparam \current_shift_inst.timer_phase.counter_10_LC_7_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_10_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_10_LC_7_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_10_LC_7_20_2  (
            .in0(N__26588),
            .in1(N__25783),
            .in2(_gnd_net_),
            .in3(N__23331),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_10 ),
            .clk(N__47337),
            .ce(N__33645),
            .sr(N__46943));
    defparam \current_shift_inst.timer_phase.counter_11_LC_7_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_11_LC_7_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_11_LC_7_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_11_LC_7_20_3  (
            .in0(N__26592),
            .in1(N__25756),
            .in2(_gnd_net_),
            .in3(N__23328),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_11 ),
            .clk(N__47337),
            .ce(N__33645),
            .sr(N__46943));
    defparam \current_shift_inst.timer_phase.counter_12_LC_7_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_12_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_12_LC_7_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_12_LC_7_20_4  (
            .in0(N__26589),
            .in1(N__26182),
            .in2(_gnd_net_),
            .in3(N__23379),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_12 ),
            .clk(N__47337),
            .ce(N__33645),
            .sr(N__46943));
    defparam \current_shift_inst.timer_phase.counter_13_LC_7_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_13_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_13_LC_7_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_13_LC_7_20_5  (
            .in0(N__26593),
            .in1(N__26152),
            .in2(_gnd_net_),
            .in3(N__23376),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_13 ),
            .clk(N__47337),
            .ce(N__33645),
            .sr(N__46943));
    defparam \current_shift_inst.timer_phase.counter_14_LC_7_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_14_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_14_LC_7_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_14_LC_7_20_6  (
            .in0(N__26590),
            .in1(N__26131),
            .in2(_gnd_net_),
            .in3(N__23373),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_14 ),
            .clk(N__47337),
            .ce(N__33645),
            .sr(N__46943));
    defparam \current_shift_inst.timer_phase.counter_15_LC_7_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_15_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_15_LC_7_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_15_LC_7_20_7  (
            .in0(N__26594),
            .in1(N__26110),
            .in2(_gnd_net_),
            .in3(N__23370),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_15 ),
            .clk(N__47337),
            .ce(N__33645),
            .sr(N__46943));
    defparam \current_shift_inst.timer_phase.counter_16_LC_7_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_16_LC_7_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_16_LC_7_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_16_LC_7_21_0  (
            .in0(N__26536),
            .in1(N__26086),
            .in2(_gnd_net_),
            .in3(N__23367),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_16 ),
            .clk(N__47331),
            .ce(N__33640),
            .sr(N__46944));
    defparam \current_shift_inst.timer_phase.counter_17_LC_7_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_17_LC_7_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_17_LC_7_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_17_LC_7_21_1  (
            .in0(N__26540),
            .in1(N__26059),
            .in2(_gnd_net_),
            .in3(N__23364),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_17 ),
            .clk(N__47331),
            .ce(N__33640),
            .sr(N__46944));
    defparam \current_shift_inst.timer_phase.counter_18_LC_7_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_18_LC_7_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_18_LC_7_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_18_LC_7_21_2  (
            .in0(N__26537),
            .in1(N__26029),
            .in2(_gnd_net_),
            .in3(N__23361),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_18 ),
            .clk(N__47331),
            .ce(N__33640),
            .sr(N__46944));
    defparam \current_shift_inst.timer_phase.counter_19_LC_7_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_19_LC_7_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_19_LC_7_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_19_LC_7_21_3  (
            .in0(N__26541),
            .in1(N__26002),
            .in2(_gnd_net_),
            .in3(N__23358),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_19 ),
            .clk(N__47331),
            .ce(N__33640),
            .sr(N__46944));
    defparam \current_shift_inst.timer_phase.counter_20_LC_7_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_20_LC_7_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_20_LC_7_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_20_LC_7_21_4  (
            .in0(N__26538),
            .in1(N__26428),
            .in2(_gnd_net_),
            .in3(N__23355),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_20 ),
            .clk(N__47331),
            .ce(N__33640),
            .sr(N__46944));
    defparam \current_shift_inst.timer_phase.counter_21_LC_7_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_21_LC_7_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_21_LC_7_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_21_LC_7_21_5  (
            .in0(N__26542),
            .in1(N__26398),
            .in2(_gnd_net_),
            .in3(N__23418),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_21 ),
            .clk(N__47331),
            .ce(N__33640),
            .sr(N__46944));
    defparam \current_shift_inst.timer_phase.counter_22_LC_7_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_22_LC_7_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_22_LC_7_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_22_LC_7_21_6  (
            .in0(N__26539),
            .in1(N__26377),
            .in2(_gnd_net_),
            .in3(N__23415),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_22 ),
            .clk(N__47331),
            .ce(N__33640),
            .sr(N__46944));
    defparam \current_shift_inst.timer_phase.counter_23_LC_7_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_23_LC_7_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_23_LC_7_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_23_LC_7_21_7  (
            .in0(N__26543),
            .in1(N__26356),
            .in2(_gnd_net_),
            .in3(N__23412),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_23 ),
            .clk(N__47331),
            .ce(N__33640),
            .sr(N__46944));
    defparam \current_shift_inst.timer_phase.counter_24_LC_7_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_24_LC_7_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_24_LC_7_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_24_LC_7_22_0  (
            .in0(N__26530),
            .in1(N__26332),
            .in2(_gnd_net_),
            .in3(N__23409),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_7_22_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_24 ),
            .clk(N__47326),
            .ce(N__33639),
            .sr(N__46946));
    defparam \current_shift_inst.timer_phase.counter_25_LC_7_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_25_LC_7_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_25_LC_7_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_25_LC_7_22_1  (
            .in0(N__26534),
            .in1(N__26305),
            .in2(_gnd_net_),
            .in3(N__23406),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_25 ),
            .clk(N__47326),
            .ce(N__33639),
            .sr(N__46946));
    defparam \current_shift_inst.timer_phase.counter_26_LC_7_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_26_LC_7_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_26_LC_7_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_26_LC_7_22_2  (
            .in0(N__26531),
            .in1(N__26257),
            .in2(_gnd_net_),
            .in3(N__23403),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_26 ),
            .clk(N__47326),
            .ce(N__33639),
            .sr(N__46946));
    defparam \current_shift_inst.timer_phase.counter_27_LC_7_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_27_LC_7_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_27_LC_7_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_27_LC_7_22_3  (
            .in0(N__26535),
            .in1(N__26212),
            .in2(_gnd_net_),
            .in3(N__23400),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_27 ),
            .clk(N__47326),
            .ce(N__33639),
            .sr(N__46946));
    defparam \current_shift_inst.timer_phase.counter_28_LC_7_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_28_LC_7_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_28_LC_7_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_28_LC_7_22_4  (
            .in0(N__26532),
            .in1(N__26279),
            .in2(_gnd_net_),
            .in3(N__23397),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_28 ),
            .clk(N__47326),
            .ce(N__33639),
            .sr(N__46946));
    defparam \current_shift_inst.timer_phase.counter_29_LC_7_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.counter_29_LC_7_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_29_LC_7_22_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_phase.counter_29_LC_7_22_5  (
            .in0(N__26234),
            .in1(N__26533),
            .in2(_gnd_net_),
            .in3(N__23394),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47326),
            .ce(N__33639),
            .sr(N__46946));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_3_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_3_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_8_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23391),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47456),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_3_7 (
            .in0(N__23562),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47456),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_6_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__23535),
            .in2(N__23553),
            .in3(N__23658),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_6_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__23520),
            .in2(N__23529),
            .in3(N__23634),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_6_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__23502),
            .in2(N__23514),
            .in3(N__23610),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_6_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__23496),
            .in2(N__23484),
            .in3(N__23586),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_6_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__23463),
            .in2(N__23475),
            .in3(N__24180),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_6_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_6_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_6_5  (
            .in0(N__24156),
            .in1(N__23442),
            .in2(N__23457),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_6_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__23424),
            .in2(N__23436),
            .in3(N__24132),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_6_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_6_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_6_7  (
            .in0(N__24108),
            .in1(N__23745),
            .in2(N__23733),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__23712),
            .in2(N__23724),
            .in3(N__24084),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__23691),
            .in2(N__23706),
            .in3(N__24015),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_8_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_8_7_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_8_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23685),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47433),
            .ce(),
            .sr(N__46850));
    defparam \pwm_generator_inst.counter_0_LC_8_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_8_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_8_8_0  (
            .in0(N__24057),
            .in1(N__23657),
            .in2(_gnd_net_),
            .in3(N__23637),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__47425),
            .ce(),
            .sr(N__46858));
    defparam \pwm_generator_inst.counter_1_LC_8_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_8_8_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_8_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_8_8_1  (
            .in0(N__24042),
            .in1(N__23633),
            .in2(_gnd_net_),
            .in3(N__23613),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__47425),
            .ce(),
            .sr(N__46858));
    defparam \pwm_generator_inst.counter_2_LC_8_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_8_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_8_8_2  (
            .in0(N__24058),
            .in1(N__23609),
            .in2(_gnd_net_),
            .in3(N__23589),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__47425),
            .ce(),
            .sr(N__46858));
    defparam \pwm_generator_inst.counter_3_LC_8_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_8_8_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_8_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_8_8_3  (
            .in0(N__24043),
            .in1(N__23585),
            .in2(_gnd_net_),
            .in3(N__23565),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__47425),
            .ce(),
            .sr(N__46858));
    defparam \pwm_generator_inst.counter_4_LC_8_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_8_8_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_8_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_8_8_4  (
            .in0(N__24059),
            .in1(N__24179),
            .in2(_gnd_net_),
            .in3(N__24159),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__47425),
            .ce(),
            .sr(N__46858));
    defparam \pwm_generator_inst.counter_5_LC_8_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_8_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_8_8_5  (
            .in0(N__24044),
            .in1(N__24154),
            .in2(_gnd_net_),
            .in3(N__24135),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__47425),
            .ce(),
            .sr(N__46858));
    defparam \pwm_generator_inst.counter_6_LC_8_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_8_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_8_8_6  (
            .in0(N__24060),
            .in1(N__24130),
            .in2(_gnd_net_),
            .in3(N__24111),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__47425),
            .ce(),
            .sr(N__46858));
    defparam \pwm_generator_inst.counter_7_LC_8_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_8_8_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_8_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_8_8_7  (
            .in0(N__24045),
            .in1(N__24107),
            .in2(_gnd_net_),
            .in3(N__24087),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__47425),
            .ce(),
            .sr(N__46858));
    defparam \pwm_generator_inst.counter_8_LC_8_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_8_9_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_8_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_8_9_0  (
            .in0(N__24047),
            .in1(N__24083),
            .in2(_gnd_net_),
            .in3(N__24063),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__47417),
            .ce(),
            .sr(N__46868));
    defparam \pwm_generator_inst.counter_9_LC_8_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_8_9_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_8_9_1  (
            .in0(N__24014),
            .in1(N__24046),
            .in2(_gnd_net_),
            .in3(N__24018),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47417),
            .ce(),
            .sr(N__46868));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_8_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_8_10_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_8_10_6  (
            .in0(N__23994),
            .in1(N__23976),
            .in2(N__23963),
            .in3(N__25122),
            .lcout(\current_shift_inst.PI_CTRL.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_8_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_8_11_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_8_11_3  (
            .in0(N__23903),
            .in1(N__23853),
            .in2(N__23823),
            .in3(N__23775),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_8_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_8_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_8_11_4  (
            .in0(N__25143),
            .in1(N__25137),
            .in2(N__25131),
            .in3(N__25128),
            .lcout(\current_shift_inst.PI_CTRL.N_47_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_8_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_8_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_8_12_1  (
            .in0(N__25733),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47392),
            .ce(N__24467),
            .sr(N__46896));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_2 .LUT_INIT=16'b1111010011000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_2  (
            .in0(N__24651),
            .in1(N__24766),
            .in2(N__25092),
            .in3(N__24969),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47392),
            .ce(N__24467),
            .sr(N__46896));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_12_5 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_8_12_5  (
            .in0(N__24970),
            .in1(N__24906),
            .in2(N__24822),
            .in3(N__24652),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47392),
            .ce(N__24467),
            .sr(N__46896));
    defparam \current_shift_inst.control_input_0_LC_8_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_8_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__26613),
            .in2(N__30708),
            .in3(N__30707),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__47382),
            .ce(N__27162),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_8_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_8_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_1_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__26604),
            .in2(_gnd_net_),
            .in3(N__24237),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__47382),
            .ce(N__27162),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_8_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_8_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__26772),
            .in2(_gnd_net_),
            .in3(N__24210),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__47382),
            .ce(N__27162),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_8_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_8_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__26754),
            .in2(_gnd_net_),
            .in3(N__24183),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__47382),
            .ce(N__27162),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_8_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_8_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_4_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__26721),
            .in2(_gnd_net_),
            .in3(N__25347),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__47382),
            .ce(N__27162),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_8_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_8_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_5_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__26688),
            .in2(_gnd_net_),
            .in3(N__25314),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__47382),
            .ce(N__27162),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_8_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_8_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_6_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__26667),
            .in2(_gnd_net_),
            .in3(N__25287),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__47382),
            .ce(N__27162),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_8_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_8_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_7_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__26658),
            .in2(_gnd_net_),
            .in3(N__25257),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__47382),
            .ce(N__27162),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_8_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_8_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_8_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__26637),
            .in2(_gnd_net_),
            .in3(N__25227),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__47376),
            .ce(N__27174),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_8_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_8_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__26946),
            .in2(_gnd_net_),
            .in3(N__25194),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__47376),
            .ce(N__27174),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_8_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_8_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_10_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__26937),
            .in2(_gnd_net_),
            .in3(N__25170),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__47376),
            .ce(N__27174),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_8_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_11_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_8_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_11_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__26928),
            .in2(_gnd_net_),
            .in3(N__25146),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_10 ),
            .carryout(\current_shift_inst.control_input_1_cry_11 ),
            .clk(N__47376),
            .ce(N__27174),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_12_LC_8_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_12_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_12_LC_8_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_12_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__26907),
            .in2(_gnd_net_),
            .in3(N__25578),
            .lcout(\current_shift_inst.control_inputZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_11 ),
            .carryout(\current_shift_inst.control_input_1_cry_12 ),
            .clk(N__47376),
            .ce(N__27174),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_13_LC_8_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_13_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_13_LC_8_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_13_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__26874),
            .in2(_gnd_net_),
            .in3(N__25554),
            .lcout(\current_shift_inst.control_inputZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_12 ),
            .carryout(\current_shift_inst.control_input_1_cry_13 ),
            .clk(N__47376),
            .ce(N__27174),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_14_LC_8_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_14_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_14_LC_8_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_14_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__26844),
            .in2(_gnd_net_),
            .in3(N__25530),
            .lcout(\current_shift_inst.control_inputZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_13 ),
            .carryout(\current_shift_inst.control_input_1_cry_14 ),
            .clk(N__47376),
            .ce(N__27174),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_15_LC_8_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_15_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_15_LC_8_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_15_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__26814),
            .in2(_gnd_net_),
            .in3(N__25506),
            .lcout(\current_shift_inst.control_inputZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_14 ),
            .carryout(\current_shift_inst.control_input_1_cry_15 ),
            .clk(N__47376),
            .ce(N__27174),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_16_LC_8_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_16_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_16_LC_8_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_16_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__26784),
            .in2(_gnd_net_),
            .in3(N__25479),
            .lcout(\current_shift_inst.control_inputZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\current_shift_inst.control_input_1_cry_16 ),
            .clk(N__47369),
            .ce(N__27184),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_17_LC_8_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_17_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_17_LC_8_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_17_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__27099),
            .in2(_gnd_net_),
            .in3(N__25452),
            .lcout(\current_shift_inst.control_inputZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_16 ),
            .carryout(\current_shift_inst.control_input_1_cry_17 ),
            .clk(N__47369),
            .ce(N__27184),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_18_LC_8_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_18_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_18_LC_8_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_18_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__27090),
            .in2(_gnd_net_),
            .in3(N__25422),
            .lcout(\current_shift_inst.control_inputZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_17 ),
            .carryout(\current_shift_inst.control_input_1_cry_18 ),
            .clk(N__47369),
            .ce(N__27184),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_19_LC_8_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_19_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_19_LC_8_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_19_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__27081),
            .in2(_gnd_net_),
            .in3(N__25395),
            .lcout(\current_shift_inst.control_inputZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_18 ),
            .carryout(\current_shift_inst.control_input_1_cry_19 ),
            .clk(N__47369),
            .ce(N__27184),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_20_LC_8_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_20_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_20_LC_8_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_20_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__27072),
            .in2(_gnd_net_),
            .in3(N__25371),
            .lcout(\current_shift_inst.control_inputZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_19 ),
            .carryout(\current_shift_inst.control_input_1_cry_20 ),
            .clk(N__47369),
            .ce(N__27184),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_21_LC_8_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_21_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_21_LC_8_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_21_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__27054),
            .in2(_gnd_net_),
            .in3(N__25713),
            .lcout(\current_shift_inst.control_inputZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_20 ),
            .carryout(\current_shift_inst.control_input_1_cry_21 ),
            .clk(N__47369),
            .ce(N__27184),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_22_LC_8_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_22_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_22_LC_8_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_22_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__27024),
            .in2(_gnd_net_),
            .in3(N__25686),
            .lcout(\current_shift_inst.control_inputZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_21 ),
            .carryout(\current_shift_inst.control_input_1_cry_22 ),
            .clk(N__47369),
            .ce(N__27184),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_23_LC_8_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_23_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_23_LC_8_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_23_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__26994),
            .in2(_gnd_net_),
            .in3(N__25659),
            .lcout(\current_shift_inst.control_inputZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_22 ),
            .carryout(\current_shift_inst.control_input_1_cry_23 ),
            .clk(N__47369),
            .ce(N__27184),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_24_LC_8_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_24_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_24_LC_8_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_24_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__26955),
            .in2(_gnd_net_),
            .in3(N__25632),
            .lcout(\current_shift_inst.control_inputZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\current_shift_inst.control_input_1_cry_24 ),
            .clk(N__47362),
            .ce(N__27186),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25629),
            .lcout(\current_shift_inst.control_input_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_8_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_8_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_8_17_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__28655),
            .in2(N__25622),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_3 ),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47355),
            .ce(N__28632),
            .sr(N__46929));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_8_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_8_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_8_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__28700),
            .in2(N__25982),
            .in3(N__25626),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47355),
            .ce(N__28632),
            .sr(N__46929));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_8_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_8_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_8_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__25955),
            .in2(N__25623),
            .in3(N__25599),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47355),
            .ce(N__28632),
            .sr(N__46929));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_8_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_8_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_8_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__25931),
            .in2(N__25983),
            .in3(N__25959),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47355),
            .ce(N__28632),
            .sr(N__46929));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_8_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_8_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_8_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__25956),
            .in2(N__25910),
            .in3(N__25935),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47355),
            .ce(N__28632),
            .sr(N__46929));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_8_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_8_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_8_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__25932),
            .in2(N__25880),
            .in3(N__25914),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47355),
            .ce(N__28632),
            .sr(N__46929));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_8_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_8_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_8_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__25851),
            .in2(N__25911),
            .in3(N__25884),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47355),
            .ce(N__28632),
            .sr(N__46929));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_8_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_8_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_8_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__25821),
            .in2(N__25881),
            .in3(N__25854),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47355),
            .ce(N__28632),
            .sr(N__46929));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_8_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_8_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_8_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__25850),
            .in2(N__25790),
            .in3(N__25824),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_11 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47346),
            .ce(N__28631),
            .sr(N__46933));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_8_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_8_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_8_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__25820),
            .in2(N__25763),
            .in3(N__25794),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47346),
            .ce(N__28631),
            .sr(N__46933));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_8_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_8_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_8_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__26189),
            .in2(N__25791),
            .in3(N__25767),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47346),
            .ce(N__28631),
            .sr(N__46933));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_8_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_8_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_8_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__26159),
            .in2(N__25764),
            .in3(N__25740),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47346),
            .ce(N__28631),
            .sr(N__46933));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_8_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_8_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_8_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__26132),
            .in2(N__26193),
            .in3(N__26166),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47346),
            .ce(N__28631),
            .sr(N__46933));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_8_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_8_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_8_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__26111),
            .in2(N__26163),
            .in3(N__26136),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47346),
            .ce(N__28631),
            .sr(N__46933));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_8_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_8_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_8_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__26133),
            .in2(N__26091),
            .in3(N__26115),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47346),
            .ce(N__28631),
            .sr(N__46933));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_8_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_8_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_8_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__26112),
            .in2(N__26064),
            .in3(N__26094),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47346),
            .ce(N__28631),
            .sr(N__46933));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_8_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_8_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__26090),
            .in2(N__26036),
            .in3(N__26067),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_19 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47338),
            .ce(N__28629),
            .sr(N__46938));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_8_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_8_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__26063),
            .in2(N__26009),
            .in3(N__26040),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47338),
            .ce(N__28629),
            .sr(N__46938));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_8_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_8_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__26435),
            .in2(N__26037),
            .in3(N__26013),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47338),
            .ce(N__28629),
            .sr(N__46938));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_8_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_8_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__26405),
            .in2(N__26010),
            .in3(N__25986),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47338),
            .ce(N__28629),
            .sr(N__46938));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_8_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_8_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__26378),
            .in2(N__26439),
            .in3(N__26412),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47338),
            .ce(N__28629),
            .sr(N__46938));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_8_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_8_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__26357),
            .in2(N__26409),
            .in3(N__26382),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47338),
            .ce(N__28629),
            .sr(N__46938));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_8_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__26379),
            .in2(N__26337),
            .in3(N__26361),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47338),
            .ce(N__28629),
            .sr(N__46938));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_8_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_8_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__26358),
            .in2(N__26310),
            .in3(N__26340),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47338),
            .ce(N__28629),
            .sr(N__46938));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_8_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_8_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__26336),
            .in2(N__26264),
            .in3(N__26313),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_27 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47332),
            .ce(N__28628),
            .sr(N__46942));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_8_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_8_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_8_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__26309),
            .in2(N__26219),
            .in3(N__26286),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47332),
            .ce(N__28628),
            .sr(N__46942));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_8_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_8_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_8_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__26283),
            .in2(N__26265),
            .in3(N__26241),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47332),
            .ce(N__28628),
            .sr(N__46942));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_8_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_8_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__26238),
            .in2(N__26220),
            .in3(N__26196),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47332),
            .ce(N__28628),
            .sr(N__46942));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_8_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_8_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_8_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26598),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47332),
            .ce(N__28628),
            .sr(N__46942));
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_8_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_8_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_8_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIB31B_LC_8_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33674),
            .lcout(\current_shift_inst.timer_phase.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_6_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_6_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_9_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26469),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47434),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_4 .LUT_INIT=16'b1000100010001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_4  (
            .in0(N__36508),
            .in1(N__37329),
            .in2(N__37869),
            .in3(N__34368),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47410),
            .ce(N__30883),
            .sr(N__46859));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_9_7 .LUT_INIT=16'b1111000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_9_9_7  (
            .in0(N__34369),
            .in1(N__37844),
            .in2(N__37366),
            .in3(N__34430),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47410),
            .ce(N__30883),
            .sr(N__46859));
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_9_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_9_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.stop_timer_s1_RNO_0_LC_9_11_5  (
            .in0(N__28982),
            .in1(N__31322),
            .in2(N__33156),
            .in3(N__31371),
            .lcout(\current_shift_inst.N_199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync0_LC_9_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync0_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync0_LC_9_12_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.S1_sync0_LC_9_12_0  (
            .in0(N__32924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.S1_syncZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47383),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_rise_LC_9_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.S1_rise_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_rise_LC_9_12_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \current_shift_inst.S1_rise_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__26445),
            .in2(_gnd_net_),
            .in3(N__26453),
            .lcout(\current_shift_inst.S1_riseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47383),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync1_LC_9_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync1_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync1_LC_9_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S1_sync1_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26460),
            .lcout(\current_shift_inst.S1_syncZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47383),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync_prev_LC_9_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync_prev_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync_prev_LC_9_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.S1_sync_prev_LC_9_12_7  (
            .in0(N__26454),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.S1_sync_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47383),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__30581),
            .in2(N__30592),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__26628),
            .in2(N__29418),
            .in3(N__30729),
            .lcout(\current_shift_inst.z_i_0_31 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__29388),
            .in2(N__28230),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_0 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__29352),
            .in2(N__28611),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_1 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__29319),
            .in2(N__26622),
            .in3(N__28671),
            .lcout(\current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_2 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__28527),
            .in2(N__28545),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_3 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__28125),
            .in2(N__28482),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_4 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__29076),
            .in2(N__28215),
            .in3(N__26607),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_5 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__28011),
            .in2(N__28005),
            .in3(N__26775),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__28170),
            .in2(N__27993),
            .in3(N__26766),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_7 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__26763),
            .in2(N__28134),
            .in3(N__26748),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_8 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__26745),
            .in2(N__26736),
            .in3(N__26715),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_9 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__26712),
            .in2(N__26703),
            .in3(N__26682),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_10 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__28236),
            .in2(N__26679),
            .in3(N__26661),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_11 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__28203),
            .in2(N__28065),
            .in3(N__26652),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_12 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__28020),
            .in2(N__26649),
            .in3(N__26631),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_13 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__28071),
            .in2(N__28386),
            .in3(N__26940),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__28119),
            .in2(N__28113),
            .in3(N__26931),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_15 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__28353),
            .in2(N__28104),
            .in3(N__26922),
            .lcout(\current_shift_inst.control_input_1_axb_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_16 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__26919),
            .in2(N__28311),
            .in3(N__26901),
            .lcout(\current_shift_inst.control_input_1_axb_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_17 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__26898),
            .in2(N__26889),
            .in3(N__26868),
            .lcout(\current_shift_inst.control_input_1_axb_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_18 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__26865),
            .in2(N__26856),
            .in3(N__26838),
            .lcout(\current_shift_inst.control_input_1_axb_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_19 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__26835),
            .in2(N__26826),
            .in3(N__26808),
            .lcout(\current_shift_inst.control_input_1_axb_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_20 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__26805),
            .in2(N__26796),
            .in3(N__26778),
            .lcout(\current_shift_inst.control_input_1_axb_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_21 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__30228),
            .in2(N__27114),
            .in3(N__27093),
            .lcout(\current_shift_inst.control_input_1_axb_17 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__30621),
            .in2(N__30609),
            .in3(N__27084),
            .lcout(\current_shift_inst.control_input_1_axb_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_23 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__30027),
            .in2(N__30744),
            .in3(N__27075),
            .lcout(\current_shift_inst.control_input_1_axb_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_24 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__30111),
            .in2(N__29151),
            .in3(N__27066),
            .lcout(\current_shift_inst.control_input_1_axb_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_25 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__27063),
            .in2(N__30369),
            .in3(N__27048),
            .lcout(\current_shift_inst.control_input_1_axb_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_26 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__27045),
            .in2(N__27036),
            .in3(N__27018),
            .lcout(\current_shift_inst.control_input_1_axb_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_27 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__27015),
            .in2(N__27006),
            .in3(N__26988),
            .lcout(\current_shift_inst.control_input_1_axb_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_28 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__26985),
            .in2(N__26973),
            .in3(N__26949),
            .lcout(\current_shift_inst.control_input_1_axb_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_29 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_25_LC_9_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_25_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_25_LC_9_17_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.control_input_25_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__30453),
            .in2(N__27255),
            .in3(N__27246),
            .lcout(\current_shift_inst.control_inputZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47347),
            .ce(N__27185),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_9_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_9_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28458),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\current_shift_inst.z_5_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_9_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_9_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__28571),
            .in2(N__27772),
            .in3(N__27135),
            .lcout(\current_shift_inst.z_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_1 ),
            .carryout(\current_shift_inst.z_5_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_9_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_9_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__27698),
            .in2(N__28589),
            .in3(N__27132),
            .lcout(\current_shift_inst.z_5_3 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_2 ),
            .carryout(\current_shift_inst.z_5_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_9_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_9_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__28493),
            .in2(N__27773),
            .in3(N__27129),
            .lcout(\current_shift_inst.z_5_4 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_3 ),
            .carryout(\current_shift_inst.z_5_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_9_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_9_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__29087),
            .in2(N__27861),
            .in3(N__27126),
            .lcout(\current_shift_inst.z_5_5 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_4 ),
            .carryout(\current_shift_inst.z_5_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_9_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_9_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__29117),
            .in2(N__27774),
            .in3(N__27123),
            .lcout(\current_shift_inst.z_5_6 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_5 ),
            .carryout(\current_shift_inst.z_5_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_9_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_9_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__27705),
            .in2(N__28187),
            .in3(N__27120),
            .lcout(\current_shift_inst.z_5_7 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_6 ),
            .carryout(\current_shift_inst.z_5_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_9_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_9_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__28147),
            .in2(N__27775),
            .in3(N__27117),
            .lcout(\current_shift_inst.z_5_8 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_7 ),
            .carryout(\current_shift_inst.z_5_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_9_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__27326),
            .in2(N__27860),
            .in3(N__27309),
            .lcout(\current_shift_inst.z_5_9 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.z_5_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_9_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__27296),
            .in2(N__27838),
            .in3(N__27279),
            .lcout(\current_shift_inst.z_5_10 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_9 ),
            .carryout(\current_shift_inst.z_5_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_9_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__28247),
            .in2(N__27857),
            .in3(N__27276),
            .lcout(\current_shift_inst.z_5_11 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_10 ),
            .carryout(\current_shift_inst.z_5_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_9_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__28280),
            .in2(N__27839),
            .in3(N__27273),
            .lcout(\current_shift_inst.z_5_12 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_11 ),
            .carryout(\current_shift_inst.z_5_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_9_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__28031),
            .in2(N__27858),
            .in3(N__27270),
            .lcout(\current_shift_inst.z_5_13 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_12 ),
            .carryout(\current_shift_inst.z_5_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_9_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__28399),
            .in2(N__27840),
            .in3(N__27267),
            .lcout(\current_shift_inst.z_5_14 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_13 ),
            .carryout(\current_shift_inst.z_5_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_9_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__28082),
            .in2(N__27859),
            .in3(N__27264),
            .lcout(\current_shift_inst.z_5_15 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_14 ),
            .carryout(\current_shift_inst.z_5_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_9_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_9_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__28364),
            .in2(N__27841),
            .in3(N__27261),
            .lcout(\current_shift_inst.z_5_16 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_15 ),
            .carryout(\current_shift_inst.z_5_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_9_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_9_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__28330),
            .in2(N__27798),
            .in3(N__27258),
            .lcout(\current_shift_inst.z_5_17 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\current_shift_inst.z_5_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_9_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_9_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__27465),
            .in2(N__27826),
            .in3(N__27441),
            .lcout(\current_shift_inst.z_5_18 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_17 ),
            .carryout(\current_shift_inst.z_5_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_9_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_9_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__27422),
            .in2(N__27799),
            .in3(N__27411),
            .lcout(\current_shift_inst.z_5_19 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_18 ),
            .carryout(\current_shift_inst.z_5_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_9_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_9_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__27395),
            .in2(N__27827),
            .in3(N__27384),
            .lcout(\current_shift_inst.z_5_20 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_19 ),
            .carryout(\current_shift_inst.z_5_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_9_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_9_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__27362),
            .in2(N__27800),
            .in3(N__27351),
            .lcout(\current_shift_inst.z_5_21 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_20 ),
            .carryout(\current_shift_inst.z_5_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_9_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_9_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__30331),
            .in2(N__27828),
            .in3(N__27348),
            .lcout(\current_shift_inst.z_5_22 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_21 ),
            .carryout(\current_shift_inst.z_5_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_9_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_9_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__30239),
            .in2(N__27801),
            .in3(N__27345),
            .lcout(\current_shift_inst.z_5_23 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_22 ),
            .carryout(\current_shift_inst.z_5_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_9_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_9_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__30664),
            .in2(N__27829),
            .in3(N__27342),
            .lcout(\current_shift_inst.z_5_24 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_23 ),
            .carryout(\current_shift_inst.z_5_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_9_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__30057),
            .in2(N__27666),
            .in3(N__27339),
            .lcout(\current_shift_inst.z_5_25 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\current_shift_inst.z_5_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_9_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__30432),
            .in2(N__27669),
            .in3(N__27948),
            .lcout(\current_shift_inst.z_5_26 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_25 ),
            .carryout(\current_shift_inst.z_5_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_9_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__27929),
            .in2(N__27667),
            .in3(N__27918),
            .lcout(\current_shift_inst.z_5_27 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_26 ),
            .carryout(\current_shift_inst.z_5_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_9_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__27902),
            .in2(N__27670),
            .in3(N__27891),
            .lcout(\current_shift_inst.z_5_28 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_27 ),
            .carryout(\current_shift_inst.z_5_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_9_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__27875),
            .in2(N__27668),
            .in3(N__27864),
            .lcout(\current_shift_inst.z_5_29 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_28 ),
            .carryout(\current_shift_inst.z_5_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_9_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__30517),
            .in2(N__27671),
            .in3(N__27489),
            .lcout(\current_shift_inst.z_5_30 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_29 ),
            .carryout(\current_shift_inst.z_5_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_9_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_9_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27486),
            .lcout(\current_shift_inst.z_5_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_10_4_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_10_4_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_10_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_10_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27483),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47435),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_10_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_10_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_10_6_7 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_10_6_7  (
            .in0(N__36752),
            .in1(N__37374),
            .in2(_gnd_net_),
            .in3(N__37698),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47418),
            .ce(N__30881),
            .sr(N__46826));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_1  (
            .in0(N__37349),
            .in1(N__37160),
            .in2(N__37242),
            .in3(N__37474),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__30885),
            .sr(N__46831));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_3  (
            .in0(N__37852),
            .in1(N__36831),
            .in2(_gnd_net_),
            .in3(N__37695),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__30885),
            .sr(N__46831));
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_10_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_10_8_0 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_22_LC_10_8_0  (
            .in0(N__41895),
            .in1(N__40800),
            .in2(N__27969),
            .in3(N__39040),
            .lcout(measured_delay_hc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47402),
            .ce(),
            .sr(N__46840));
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_10_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_10_8_6 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_20_LC_10_8_6  (
            .in0(N__28958),
            .in1(N__40799),
            .in2(N__41901),
            .in3(N__39039),
            .lcout(measured_delay_hc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47402),
            .ce(),
            .sr(N__46840));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_5_LC_10_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_5_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_5_LC_10_9_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_5_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__36562),
            .in2(_gnd_net_),
            .in3(N__37038),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_10_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_10_9_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_10_9_1  (
            .in0(N__27964),
            .in1(N__28897),
            .in2(N__27984),
            .in3(N__31212),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto31_LC_10_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto31_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto31_LC_10_9_2 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto31_LC_10_9_2  (
            .in0(N__37842),
            .in1(N__29028),
            .in2(N__27981),
            .in3(N__29052),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_9_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_9_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_10_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27978),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47393),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_10_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_10_9_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_10_9_4  (
            .in0(N__28898),
            .in1(N__27965),
            .in2(N__28959),
            .in3(N__29051),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_c_LC_10_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_c_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_c_LC_10_9_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto31_c_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27951),
            .in3(N__37843),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto31_cZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_10_10_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_10_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_10_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_11_LC_10_10_6  (
            .in0(N__37485),
            .in1(N__36655),
            .in2(N__37367),
            .in3(N__37141),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47384),
            .ce(N__37107),
            .sr(N__46851));
    defparam \current_shift_inst.meas_state_0_LC_10_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.meas_state_0_LC_10_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.meas_state_0_LC_10_11_0 .LUT_INIT=16'b0111111110101010;
    LogicCell40 \current_shift_inst.meas_state_0_LC_10_11_0  (
            .in0(N__31373),
            .in1(N__28987),
            .in2(N__33155),
            .in3(N__31334),
            .lcout(\current_shift_inst.meas_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47377),
            .ce(),
            .sr(N__46860));
    defparam \current_shift_inst.phase_valid_LC_10_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.phase_valid_LC_10_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.phase_valid_LC_10_11_1 .LUT_INIT=16'b1010100011111000;
    LogicCell40 \current_shift_inst.phase_valid_LC_10_11_1  (
            .in0(N__31333),
            .in1(N__31425),
            .in2(N__28994),
            .in3(N__31372),
            .lcout(\current_shift_inst.phase_validZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47377),
            .ce(),
            .sr(N__46860));
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_10_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_10_11_6 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_23_LC_10_11_6  (
            .in0(N__29067),
            .in1(N__40801),
            .in2(N__41852),
            .in3(N__39037),
            .lcout(measured_delay_hc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47377),
            .ce(),
            .sr(N__46860));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_10_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_10_12_0 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_10_12_0  (
            .in0(N__29522),
            .in1(N__28049),
            .in2(N__29571),
            .in3(N__28302),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_10_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_10_12_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28053),
            .in3(N__29521),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_10_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_10_12_7 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_27_LC_10_12_7  (
            .in0(N__29172),
            .in1(N__40802),
            .in2(N__41900),
            .in3(N__39038),
            .lcout(measured_delay_hc_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47371),
            .ce(),
            .sr(N__46872));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_13_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_13_0  (
            .in0(N__29217),
            .in1(N__28195),
            .in2(N__29136),
            .in3(N__29759),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__29132),
            .in2(_gnd_net_),
            .in3(N__29216),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_13_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__28196),
            .in2(_gnd_net_),
            .in3(N__29758),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__29101),
            .in2(_gnd_net_),
            .in3(N__29249),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__28300),
            .in2(_gnd_net_),
            .in3(N__29567),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_13_5 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_13_5  (
            .in0(N__28197),
            .in1(N__28160),
            .in2(N__29717),
            .in3(N__29760),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28164),
            .in3(N__29710),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7  (
            .in0(N__28515),
            .in1(N__29248),
            .in2(N__29292),
            .in3(N__29102),
            .lcout(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0  (
            .in0(N__28095),
            .in1(N__28375),
            .in2(N__30015),
            .in3(N__29978),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__28094),
            .in2(_gnd_net_),
            .in3(N__30010),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI190J_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__28376),
            .in2(_gnd_net_),
            .in3(N__29977),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3  (
            .in0(N__28416),
            .in1(N__28093),
            .in2(N__29487),
            .in3(N__30011),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_14_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__28415),
            .in2(_gnd_net_),
            .in3(N__29483),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_14_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_14_5  (
            .in0(N__28377),
            .in1(N__28346),
            .in2(N__29982),
            .in3(N__29942),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__29941),
            .in2(_gnd_net_),
            .in3(N__28347),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_10_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_10_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_10_14_7  (
            .in0(N__29606),
            .in1(N__28301),
            .in2(N__28269),
            .in3(N__29563),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_10_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_10_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_10_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31869),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47349),
            .ce(N__31694),
            .sr(N__46900));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31836),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47349),
            .ce(N__31694),
            .sr(N__46900));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31673),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47349),
            .ce(N__31694),
            .sr(N__46900));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_15_3  (
            .in0(N__31674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47349),
            .ce(N__31694),
            .sr(N__46900));
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_16_0 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_16_0  (
            .in0(N__30560),
            .in1(N__28451),
            .in2(_gnd_net_),
            .in3(N__29384),
            .lcout(\current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_10_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_10_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_10_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28701),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47340),
            .ce(N__28630),
            .sr(N__46908));
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_10_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_10_16_2 .LUT_INIT=16'b0101010101100101;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_10_16_2  (
            .in0(N__28595),
            .in1(N__28566),
            .in2(N__30579),
            .in3(N__28450),
            .lcout(\current_shift_inst.N_1633_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_10_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_10_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_10_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28659),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47340),
            .ce(N__28630),
            .sr(N__46908));
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_16_4 .LUT_INIT=16'b1001101010011010;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_16_4  (
            .in0(N__28570),
            .in1(N__28452),
            .in2(N__30580),
            .in3(N__29348),
            .lcout(\current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_10_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_10_16_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_10_16_5  (
            .in0(N__28453),
            .in1(N__28596),
            .in2(N__28572),
            .in3(N__30564),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ),
            .ltout(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__28507),
            .in2(N__28530),
            .in3(N__29280),
            .lcout(\current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_16_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_16_7  (
            .in0(N__29281),
            .in1(_gnd_net_),
            .in2(N__28514),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_17_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_17_0  (
            .in0(N__29442),
            .in1(N__29408),
            .in2(N__28467),
            .in3(_gnd_net_),
            .lcout(G_406),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\current_shift_inst.z_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__29380),
            .in2(N__28425),
            .in3(N__28457),
            .lcout(G_405),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_0 ),
            .carryout(\current_shift_inst.z_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__29344),
            .in2(N__28764),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_1 ),
            .carryout(\current_shift_inst.z_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__29312),
            .in2(N__28755),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_2 ),
            .carryout(\current_shift_inst.z_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__28746),
            .in2(N__29285),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_3 ),
            .carryout(\current_shift_inst.z_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__29239),
            .in2(N__28740),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_4 ),
            .carryout(\current_shift_inst.z_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__29203),
            .in2(N__28731),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_5 ),
            .carryout(\current_shift_inst.z_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__28722),
            .in2(N__29749),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_6 ),
            .carryout(\current_shift_inst.z_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__28716),
            .in2(N__29701),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\current_shift_inst.z_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__28707),
            .in2(N__29659),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_8 ),
            .carryout(\current_shift_inst.z_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__28821),
            .in2(N__29627),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_9 ),
            .carryout(\current_shift_inst.z_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__28815),
            .in2(N__29593),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_10 ),
            .carryout(\current_shift_inst.z_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(N__28809),
            .in2(N__29559),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_11 ),
            .carryout(\current_shift_inst.z_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__28803),
            .in2(N__29512),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_12 ),
            .carryout(\current_shift_inst.z_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__28797),
            .in2(N__29473),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_13 ),
            .carryout(\current_shift_inst.z_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__28791),
            .in2(N__30002),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_14 ),
            .carryout(\current_shift_inst.z_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__28785),
            .in2(N__29969),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\current_shift_inst.z_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__28776),
            .in2(N__29931),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_16 ),
            .carryout(\current_shift_inst.z_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__28770),
            .in2(N__29893),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_17 ),
            .carryout(\current_shift_inst.z_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__28875),
            .in2(N__29852),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_18 ),
            .carryout(\current_shift_inst.z_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__29819),
            .in2(N__28869),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_19 ),
            .carryout(\current_shift_inst.z_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__28860),
            .in2(N__29792),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_20 ),
            .carryout(\current_shift_inst.z_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__28854),
            .in2(N__30280),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_21 ),
            .carryout(\current_shift_inst.z_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__28848),
            .in2(N__30312),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_22 ),
            .carryout(\current_shift_inst.z_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__28842),
            .in2(N__30647),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\current_shift_inst.z_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__30093),
            .in2(N__28836),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_24 ),
            .carryout(\current_shift_inst.z_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__28827),
            .in2(N__30398),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_25 ),
            .carryout(\current_shift_inst.z_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__28938),
            .in2(N__30188),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_26 ),
            .carryout(\current_shift_inst.z_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__28932),
            .in2(N__30158),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_27 ),
            .carryout(\current_shift_inst.z_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__30128),
            .in2(N__28926),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_28 ),
            .carryout(\current_shift_inst.z_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__30469),
            .in2(N__28917),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_29 ),
            .carryout(\current_shift_inst.z_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_10_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_10_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.un10_control_input_z_s_31_LC_10_20_7  (
            .in0(N__30593),
            .in1(N__28908),
            .in2(N__30500),
            .in3(N__28902),
            .lcout(\current_shift_inst.z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_11_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_11_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_11_5_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_11_5_5  (
            .in0(N__37848),
            .in1(N__37751),
            .in2(_gnd_net_),
            .in3(N__37689),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47419),
            .ce(N__30887),
            .sr(N__46816));
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_11_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_11_6_5 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_21_LC_11_6_5  (
            .in0(N__41880),
            .in1(N__40759),
            .in2(N__28899),
            .in3(N__39042),
            .lcout(measured_delay_hc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47412),
            .ce(),
            .sr(N__46821));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_d_LC_11_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_d_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_d_LC_11_7_2 .LUT_INIT=16'b1111001111110111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto31_d_LC_11_7_2  (
            .in0(N__40554),
            .in1(N__31191),
            .in2(N__37870),
            .in3(N__31443),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0 ),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto31_dZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_11_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_11_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_11_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_0_LC_11_7_3  (
            .in0(N__37361),
            .in1(N__37161),
            .in2(N__28878),
            .in3(N__36992),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(N__30882),
            .sr(N__46827));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_11_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_11_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_11_7_6  (
            .in0(N__37162),
            .in1(N__36606),
            .in2(N__37409),
            .in3(N__37469),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(N__30882),
            .sr(N__46827));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_0  (
            .in0(N__37471),
            .in1(N__37323),
            .in2(N__36660),
            .in3(N__37155),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47394),
            .ce(N__30856),
            .sr(N__46832));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_11_8_1  (
            .in0(N__37322),
            .in1(N__37154),
            .in2(N__40563),
            .in3(N__37473),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47394),
            .ce(N__30856),
            .sr(N__46832));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_11_8_2  (
            .in0(N__37472),
            .in1(N__37324),
            .in2(N__37566),
            .in3(N__37156),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47394),
            .ce(N__30856),
            .sr(N__46832));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_3  (
            .in0(N__36702),
            .in1(N__37153),
            .in2(N__37365),
            .in3(N__37470),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47394),
            .ce(N__30856),
            .sr(N__46832));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_8_4 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_11_8_4  (
            .in0(N__37651),
            .in1(N__36792),
            .in2(_gnd_net_),
            .in3(N__37328),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47394),
            .ce(N__30856),
            .sr(N__46832));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_5  (
            .in0(N__37321),
            .in1(N__37047),
            .in2(_gnd_net_),
            .in3(N__37652),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47394),
            .ce(N__30856),
            .sr(N__46832));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_9_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_9_1  (
            .in0(N__36230),
            .in1(N__32735),
            .in2(_gnd_net_),
            .in3(N__32813),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_9_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_9_4  (
            .in0(N__28954),
            .in1(N__40541),
            .in2(_gnd_net_),
            .in3(N__36827),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_9_5  (
            .in0(N__36563),
            .in1(N__36791),
            .in2(N__36512),
            .in3(N__34422),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_3_LC_11_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_3_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_3_LC_11_10_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_14_3_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__32949),
            .in2(_gnd_net_),
            .in3(N__29066),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_LC_11_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_LC_11_10_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_14_LC_11_10_1  (
            .in0(N__32966),
            .in1(N__32895),
            .in2(N__29055),
            .in3(N__29160),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_11_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_11_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_11_10_2  (
            .in0(N__36784),
            .in1(N__36751),
            .in2(N__36516),
            .in3(N__37561),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_11_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_11_10_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_11_10_5  (
            .in0(N__36241),
            .in1(N__32803),
            .in2(_gnd_net_),
            .in3(N__32760),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto3_LC_11_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto3_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto3_LC_11_10_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto3_LC_11_10_6  (
            .in0(N__36875),
            .in1(N__36915),
            .in2(_gnd_net_),
            .in3(N__40886),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlt30_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_6_LC_11_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_6_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_6_LC_11_10_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_14_6_LC_11_10_7  (
            .in0(N__29043),
            .in1(N__31203),
            .in2(N__29037),
            .in3(N__29034),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_11_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_11_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__33370),
            .in2(_gnd_net_),
            .in3(N__33114),
            .lcout(\current_shift_inst.timer_s1.N_187_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.start_timer_s1_LC_11_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.start_timer_s1_LC_11_11_3 .LUT_INIT=16'b0100111111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_11_11_3  (
            .in0(N__28986),
            .in1(N__33141),
            .in2(N__31344),
            .in3(N__31392),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47372),
            .ce(N__34786),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_11_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_11_4  (
            .in0(N__33140),
            .in1(N__33371),
            .in2(_gnd_net_),
            .in3(N__33115),
            .lcout(\current_shift_inst.timer_s1.N_191_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_phase_LC_11_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_phase_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.stop_timer_phase_LC_11_11_6 .LUT_INIT=16'b1101110111000000;
    LogicCell40 \current_shift_inst.stop_timer_phase_LC_11_11_6  (
            .in0(N__31393),
            .in1(N__31342),
            .in2(N__31421),
            .in3(N__33729),
            .lcout(\current_shift_inst.stop_timer_phaseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47372),
            .ce(N__34786),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_12_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_11_12_0  (
            .in0(N__33095),
            .in1(N__33068),
            .in2(N__46988),
            .in3(N__34291),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47364),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_11_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_11_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_11_12_6  (
            .in0(N__31286),
            .in1(N__31301),
            .in2(N__31275),
            .in3(N__29171),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__30072),
            .in2(_gnd_net_),
            .in3(N__30099),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_11_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_11_13_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_11_13_2  (
            .in0(N__29250),
            .in1(N__29131),
            .in2(N__29106),
            .in3(N__29210),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_11_14_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_11_14_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_0_LC_11_14_0  (
            .in0(N__45673),
            .in1(N__45379),
            .in2(N__45599),
            .in3(N__41089),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(N__34793),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_11_14_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_11_14_1 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_1_LC_11_14_1  (
            .in0(N__41090),
            .in1(N__45590),
            .in2(N__45413),
            .in3(N__45674),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(N__34793),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_0_LC_11_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_11_14_2 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_11_14_2  (
            .in0(N__36302),
            .in1(N__35119),
            .in2(_gnd_net_),
            .in3(N__35106),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(N__34793),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_state_0_LC_11_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_11_14_4 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_11_14_4  (
            .in0(N__33096),
            .in1(N__33061),
            .in2(_gnd_net_),
            .in3(N__34293),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(N__34793),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29184),
            .lcout(\current_shift_inst.un4_control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29178),
            .lcout(\current_shift_inst.un4_control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_14_7  (
            .in0(N__31260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_11_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_11_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_11_15_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_11_15_0  (
            .in0(N__37697),
            .in1(N__37885),
            .in2(_gnd_net_),
            .in3(N__37941),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47341),
            .ce(N__30886),
            .sr(N__46887));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_15_1 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_11_15_1  (
            .in0(N__37884),
            .in1(N__36564),
            .in2(_gnd_net_),
            .in3(N__37696),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47341),
            .ce(N__30886),
            .sr(N__46887));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_15_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__31503),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31494),
            .lcout(\current_shift_inst.un4_control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31485),
            .lcout(\current_shift_inst.un4_control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31476),
            .lcout(\current_shift_inst.un4_control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31467),
            .lcout(\current_shift_inst.un4_control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31458),
            .lcout(\current_shift_inst.un4_control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__29451),
            .in2(N__29441),
            .in3(N__29440),
            .lcout(\current_shift_inst.un38_control_input_0 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__29397),
            .in2(_gnd_net_),
            .in3(N__29364),
            .lcout(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__29361),
            .in2(_gnd_net_),
            .in3(N__29328),
            .lcout(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__29325),
            .in2(_gnd_net_),
            .in3(N__29301),
            .lcout(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__29298),
            .in2(_gnd_net_),
            .in3(N__29259),
            .lcout(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__29256),
            .in2(_gnd_net_),
            .in3(N__29226),
            .lcout(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__29223),
            .in2(_gnd_net_),
            .in3(N__29187),
            .lcout(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__29766),
            .in2(_gnd_net_),
            .in3(N__29730),
            .lcout(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__29727),
            .in2(_gnd_net_),
            .in3(N__29676),
            .lcout(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__33186),
            .in2(_gnd_net_),
            .in3(N__29640),
            .lcout(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__33168),
            .in2(_gnd_net_),
            .in3(N__29610),
            .lcout(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__33504),
            .in2(_gnd_net_),
            .in3(N__29574),
            .lcout(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__33468),
            .in2(_gnd_net_),
            .in3(N__29532),
            .lcout(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__33450),
            .in2(_gnd_net_),
            .in3(N__29490),
            .lcout(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__33420),
            .in2(_gnd_net_),
            .in3(N__29454),
            .lcout(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__33402),
            .in2(_gnd_net_),
            .in3(N__29985),
            .lcout(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__33384),
            .in2(_gnd_net_),
            .in3(N__29952),
            .lcout(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__33486),
            .in2(_gnd_net_),
            .in3(N__29910),
            .lcout(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_18_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31593),
            .in3(N__29868),
            .lcout(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__31623),
            .in2(_gnd_net_),
            .in3(N__29835),
            .lcout(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__33204),
            .in2(_gnd_net_),
            .in3(N__29808),
            .lcout(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__31875),
            .in2(_gnd_net_),
            .in3(N__29775),
            .lcout(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__33432),
            .in2(_gnd_net_),
            .in3(N__29772),
            .lcout(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__32985),
            .in2(_gnd_net_),
            .in3(N__29769),
            .lcout(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__31890),
            .in2(_gnd_net_),
            .in3(N__30213),
            .lcout(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__31575),
            .in2(_gnd_net_),
            .in3(N__30210),
            .lcout(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__31563),
            .in2(_gnd_net_),
            .in3(N__30207),
            .lcout(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__31638),
            .in2(_gnd_net_),
            .in3(N__30171),
            .lcout(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__31653),
            .in2(_gnd_net_),
            .in3(N__30141),
            .lcout(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_19_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31611),
            .in3(N__30117),
            .lcout(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_29 ),
            .carryout(\current_shift_inst.un4_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_19_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_19_6  (
            .in0(N__30585),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30114),
            .lcout(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_11_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_11_19_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_11_19_7  (
            .in0(N__30098),
            .in1(N__30439),
            .in2(N__30071),
            .in3(N__30394),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_20_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_20_0  (
            .in0(N__30646),
            .in1(N__30094),
            .in2(N__30684),
            .in3(N__30070),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_20_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_20_1  (
            .in0(N__30645),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30679),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_11_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_11_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_i_31_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30722),
            .lcout(\current_shift_inst.z_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_20_3 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_20_3  (
            .in0(N__30683),
            .in1(N__30315),
            .in2(N__30648),
            .in3(N__30254),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_4  (
            .in0(N__30314),
            .in1(_gnd_net_),
            .in2(N__30255),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_0_25_LC_11_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_11_20_5 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \current_shift_inst.control_input_RNO_0_25_LC_11_20_5  (
            .in0(N__30594),
            .in1(N__30525),
            .in2(N__30501),
            .in3(N__30473),
            .lcout(\current_shift_inst.un38_control_input_0_axb_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__30440),
            .in2(_gnd_net_),
            .in3(N__30393),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_11_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_11_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_11_20_7  (
            .in0(N__30350),
            .in1(N__30313),
            .in2(N__30291),
            .in3(N__30250),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_LC_11_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_LC_11_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.running_LC_11_22_7 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_phase.running_LC_11_22_7  (
            .in0(N__33705),
            .in1(N__33673),
            .in2(_gnd_net_),
            .in3(N__33743),
            .lcout(\current_shift_inst.timer_phase.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47310),
            .ce(),
            .sr(N__46934));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_3_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_3_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_12_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30900),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47426),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_12_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_12_5_6 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_12_5_6  (
            .in0(N__37936),
            .in1(N__37234),
            .in2(_gnd_net_),
            .in3(N__37046),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_5_7 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_5_7  (
            .in0(N__36753),
            .in1(N__34305),
            .in2(N__30891),
            .in3(N__34323),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_12_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_12_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_12_6_0 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_12_6_0  (
            .in0(N__37668),
            .in1(N__36871),
            .in2(_gnd_net_),
            .in3(N__37373),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47401),
            .ce(N__30884),
            .sr(N__46817));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_12_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_12_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_12_6_2 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_12_6_2  (
            .in0(N__37667),
            .in1(N__37372),
            .in2(_gnd_net_),
            .in3(N__36913),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47401),
            .ce(N__30884),
            .sr(N__46817));
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_12_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_12_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_12_6_5 .LUT_INIT=16'b1010000010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_12_6_5  (
            .in0(N__37371),
            .in1(_gnd_net_),
            .in2(N__36955),
            .in3(N__37666),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47401),
            .ce(N__30884),
            .sr(N__46817));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_12_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_12_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__30795),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__30774),
            .in2(N__30786),
            .in3(N__33820),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__30750),
            .in2(N__30768),
            .in3(N__33803),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__31038),
            .in2(N__31050),
            .in3(N__33767),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__31020),
            .in2(N__31032),
            .in3(N__34070),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__30999),
            .in2(N__31014),
            .in3(N__34049),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(N__30978),
            .in2(N__30993),
            .in3(N__34028),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__30960),
            .in2(N__30972),
            .in3(N__34004),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__30939),
            .in2(N__30954),
            .in3(N__33980),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__30924),
            .in2(N__30933),
            .in3(N__33953),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_8_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_8_2  (
            .in0(N__33932),
            .in1(N__30906),
            .in2(N__30918),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__31161),
            .in2(N__31173),
            .in3(N__34253),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__31146),
            .in2(N__31155),
            .in3(N__34229),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__31128),
            .in2(N__31140),
            .in3(N__34208),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__31107),
            .in2(N__31122),
            .in3(N__34187),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__31089),
            .in2(N__31101),
            .in3(N__34166),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__31074),
            .in2(N__31083),
            .in3(N__34143),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_9_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_9_1  (
            .in0(N__34115),
            .in1(N__31056),
            .in2(N__31068),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__31242),
            .in2(N__31254),
            .in3(N__34094),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__31221),
            .in2(N__31236),
            .in3(N__34346),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31215),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_9_6  (
            .in0(N__37223),
            .in1(N__36609),
            .in2(N__37940),
            .in3(N__36656),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_12_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_12_9_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_12_9_7  (
            .in0(N__34634),
            .in1(N__33824),
            .in2(_gnd_net_),
            .in3(N__34582),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_12_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_12_10_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__32796),
            .in2(_gnd_net_),
            .in3(N__32682),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_10_2  (
            .in0(N__36951),
            .in1(N__36701),
            .in2(N__34431),
            .in3(N__37752),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync_prev_LC_12_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync_prev_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync_prev_LC_12_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S3_sync_prev_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33012),
            .lcout(\current_shift_inst.S3_sync_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47370),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_rise_LC_12_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.S3_rise_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_rise_LC_12_10_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \current_shift_inst.S3_rise_LC_12_10_6  (
            .in0(N__33011),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31197),
            .lcout(\current_shift_inst.S3_riseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47370),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_3_LC_12_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_3_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_3_LC_12_10_7 .LUT_INIT=16'b0000110001001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_3_LC_12_10_7  (
            .in0(N__40555),
            .in1(N__34381),
            .in2(N__31190),
            .in3(N__31442),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.start_timer_phase_LC_12_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_phase_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.start_timer_phase_LC_12_11_3 .LUT_INIT=16'b0101110101001100;
    LogicCell40 \current_shift_inst.start_timer_phase_LC_12_11_3  (
            .in0(N__31335),
            .in1(N__33689),
            .in2(N__31420),
            .in3(N__31394),
            .lcout(\current_shift_inst.start_timer_phaseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47363),
            .ce(N__34785),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_12_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_12_11_6 .LUT_INIT=16'b0100000001100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_12_11_6  (
            .in0(N__32750),
            .in1(N__32812),
            .in2(N__36246),
            .in3(N__34589),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47363),
            .ce(N__34785),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_LC_12_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.stop_timer_s1_LC_12_11_7 .LUT_INIT=16'b1111110111001100;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_12_11_7  (
            .in0(N__31395),
            .in1(N__31353),
            .in2(N__31343),
            .in3(N__33117),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47363),
            .ce(N__34785),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.prev_hc_sig_LC_12_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_hc_sig_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_hc_sig_LC_12_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.prev_hc_sig_LC_12_12_1  (
            .in0(N__34292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.prev_hc_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47356),
            .ce(),
            .sr(N__46852));
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_12_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_12_12_3 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_28_LC_12_12_3  (
            .in0(N__31302),
            .in1(N__40834),
            .in2(N__41892),
            .in3(N__39027),
            .lcout(measured_delay_hc_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47356),
            .ce(),
            .sr(N__46852));
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_12_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_12_12_4 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_29_LC_12_12_4  (
            .in0(N__39028),
            .in1(N__41869),
            .in2(N__31290),
            .in3(N__40836),
            .lcout(measured_delay_hc_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47356),
            .ce(),
            .sr(N__46852));
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_12_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_12_12_5 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_30_LC_12_12_5  (
            .in0(N__31274),
            .in1(N__40835),
            .in2(N__41893),
            .in3(N__39029),
            .lcout(measured_delay_hc_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47356),
            .ce(),
            .sr(N__46852));
    defparam \phase_controller_inst1.T01_er_LC_12_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_er_LC_12_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_er_LC_12_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.T01_er_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34458),
            .lcout(shift_flag_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47348),
            .ce(N__33024),
            .sr(N__46861));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_14_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__31802),
            .in2(N__31868),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47339),
            .ce(N__31698),
            .sr(N__46873));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__31781),
            .in2(N__31835),
            .in3(N__31497),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47339),
            .ce(N__31698),
            .sr(N__46873));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__31803),
            .in2(N__31761),
            .in3(N__31488),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47339),
            .ce(N__31698),
            .sr(N__46873));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__31782),
            .in2(N__31731),
            .in3(N__31479),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47339),
            .ce(N__31698),
            .sr(N__46873));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__31757),
            .in2(N__32138),
            .in3(N__31470),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47339),
            .ce(N__31698),
            .sr(N__46873));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__31727),
            .in2(N__32111),
            .in3(N__31461),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47339),
            .ce(N__31698),
            .sr(N__46873));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__32081),
            .in2(N__32139),
            .in3(N__31452),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47339),
            .ce(N__31698),
            .sr(N__46873));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__32054),
            .in2(N__32112),
            .in3(N__31449),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47339),
            .ce(N__31698),
            .sr(N__46873));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__32082),
            .in2(N__32030),
            .in3(N__31446),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47333),
            .ce(N__31697),
            .sr(N__46881));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__32055),
            .in2(N__32003),
            .in3(N__31530),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47333),
            .ce(N__31697),
            .sr(N__46881));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__31976),
            .in2(N__32031),
            .in3(N__31527),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47333),
            .ce(N__31697),
            .sr(N__46881));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__31955),
            .in2(N__32004),
            .in3(N__31524),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47333),
            .ce(N__31697),
            .sr(N__46881));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__31977),
            .in2(N__31932),
            .in3(N__31521),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47333),
            .ce(N__31697),
            .sr(N__46881));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__31956),
            .in2(N__32357),
            .in3(N__31518),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47333),
            .ce(N__31697),
            .sr(N__46881));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__31928),
            .in2(N__32328),
            .in3(N__31515),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47333),
            .ce(N__31697),
            .sr(N__46881));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__32297),
            .in2(N__32358),
            .in3(N__31512),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47333),
            .ce(N__31697),
            .sr(N__46881));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__32327),
            .in2(N__32270),
            .in3(N__31509),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47327),
            .ce(N__31696),
            .sr(N__46888));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__32298),
            .in2(N__32240),
            .in3(N__31506),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47327),
            .ce(N__31696),
            .sr(N__46888));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__32210),
            .in2(N__32271),
            .in3(N__31557),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47327),
            .ce(N__31696),
            .sr(N__46888));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__32186),
            .in2(N__32241),
            .in3(N__31554),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47327),
            .ce(N__31696),
            .sr(N__46888));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__32211),
            .in2(N__32165),
            .in3(N__31551),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47327),
            .ce(N__31696),
            .sr(N__46888));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__32187),
            .in2(N__32591),
            .in3(N__31548),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47327),
            .ce(N__31696),
            .sr(N__46888));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__32561),
            .in2(N__32166),
            .in3(N__31545),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47327),
            .ce(N__31696),
            .sr(N__46888));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__32531),
            .in2(N__32592),
            .in3(N__31542),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47327),
            .ce(N__31696),
            .sr(N__46888));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__32562),
            .in2(N__32504),
            .in3(N__31539),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47322),
            .ce(N__31695),
            .sr(N__46901));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__32474),
            .in2(N__32535),
            .in3(N__31536),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47322),
            .ce(N__31695),
            .sr(N__46901));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__32454),
            .in2(N__32505),
            .in3(N__31533),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47322),
            .ce(N__31695),
            .sr(N__46901));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__32475),
            .in2(N__32430),
            .in3(N__31701),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47322),
            .ce(N__31695),
            .sr(N__46901));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31677),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31659),
            .lcout(\current_shift_inst.un4_control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_18_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__31644),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31632),
            .lcout(\current_shift_inst.un4_control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31617),
            .lcout(\current_shift_inst.un4_control_input_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_18_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__31602),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31584),
            .lcout(\current_shift_inst.un4_control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_18_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_18_5  (
            .in0(N__31569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31899),
            .lcout(\current_shift_inst.un4_control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_18_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_18_7  (
            .in0(N__31884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_12_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_12_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_12_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_12_19_0  (
            .in0(N__33315),
            .in1(N__31858),
            .in2(_gnd_net_),
            .in3(N__31839),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__47315),
            .ce(N__32403),
            .sr(N__46914));
    defparam \current_shift_inst.timer_s1.counter_1_LC_12_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_12_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_12_19_1  (
            .in0(N__33307),
            .in1(N__31825),
            .in2(_gnd_net_),
            .in3(N__31806),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__47315),
            .ce(N__32403),
            .sr(N__46914));
    defparam \current_shift_inst.timer_s1.counter_2_LC_12_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_12_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_12_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_12_19_2  (
            .in0(N__33316),
            .in1(N__31801),
            .in2(_gnd_net_),
            .in3(N__31785),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__47315),
            .ce(N__32403),
            .sr(N__46914));
    defparam \current_shift_inst.timer_s1.counter_3_LC_12_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_12_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_12_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_12_19_3  (
            .in0(N__33308),
            .in1(N__31780),
            .in2(_gnd_net_),
            .in3(N__31764),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__47315),
            .ce(N__32403),
            .sr(N__46914));
    defparam \current_shift_inst.timer_s1.counter_4_LC_12_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_12_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_12_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_12_19_4  (
            .in0(N__33317),
            .in1(N__31753),
            .in2(_gnd_net_),
            .in3(N__31734),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__47315),
            .ce(N__32403),
            .sr(N__46914));
    defparam \current_shift_inst.timer_s1.counter_5_LC_12_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_12_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_12_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_12_19_5  (
            .in0(N__33309),
            .in1(N__31723),
            .in2(_gnd_net_),
            .in3(N__31704),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__47315),
            .ce(N__32403),
            .sr(N__46914));
    defparam \current_shift_inst.timer_s1.counter_6_LC_12_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_12_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_12_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_12_19_6  (
            .in0(N__33318),
            .in1(N__32131),
            .in2(_gnd_net_),
            .in3(N__32115),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__47315),
            .ce(N__32403),
            .sr(N__46914));
    defparam \current_shift_inst.timer_s1.counter_7_LC_12_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_12_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_12_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_12_19_7  (
            .in0(N__33310),
            .in1(N__32099),
            .in2(_gnd_net_),
            .in3(N__32085),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__47315),
            .ce(N__32403),
            .sr(N__46914));
    defparam \current_shift_inst.timer_s1.counter_8_LC_12_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_12_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_12_20_0  (
            .in0(N__33335),
            .in1(N__32074),
            .in2(_gnd_net_),
            .in3(N__32058),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__47312),
            .ce(N__32411),
            .sr(N__46921));
    defparam \current_shift_inst.timer_s1.counter_9_LC_12_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_12_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_12_20_1  (
            .in0(N__33322),
            .in1(N__32053),
            .in2(_gnd_net_),
            .in3(N__32034),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__47312),
            .ce(N__32411),
            .sr(N__46921));
    defparam \current_shift_inst.timer_s1.counter_10_LC_12_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_12_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_12_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_12_20_2  (
            .in0(N__33332),
            .in1(N__32023),
            .in2(_gnd_net_),
            .in3(N__32007),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__47312),
            .ce(N__32411),
            .sr(N__46921));
    defparam \current_shift_inst.timer_s1.counter_11_LC_12_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_12_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_12_20_3  (
            .in0(N__33319),
            .in1(N__31996),
            .in2(_gnd_net_),
            .in3(N__31980),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__47312),
            .ce(N__32411),
            .sr(N__46921));
    defparam \current_shift_inst.timer_s1.counter_12_LC_12_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_12_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_12_20_4  (
            .in0(N__33333),
            .in1(N__31975),
            .in2(_gnd_net_),
            .in3(N__31959),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__47312),
            .ce(N__32411),
            .sr(N__46921));
    defparam \current_shift_inst.timer_s1.counter_13_LC_12_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_12_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_12_20_5  (
            .in0(N__33320),
            .in1(N__31949),
            .in2(_gnd_net_),
            .in3(N__31935),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__47312),
            .ce(N__32411),
            .sr(N__46921));
    defparam \current_shift_inst.timer_s1.counter_14_LC_12_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_12_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_12_20_6  (
            .in0(N__33334),
            .in1(N__31924),
            .in2(_gnd_net_),
            .in3(N__31902),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__47312),
            .ce(N__32411),
            .sr(N__46921));
    defparam \current_shift_inst.timer_s1.counter_15_LC_12_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_12_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_12_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_12_20_7  (
            .in0(N__33321),
            .in1(N__32345),
            .in2(_gnd_net_),
            .in3(N__32331),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__47312),
            .ce(N__32411),
            .sr(N__46921));
    defparam \current_shift_inst.timer_s1.counter_16_LC_12_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_12_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_12_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_12_21_0  (
            .in0(N__33311),
            .in1(N__32317),
            .in2(_gnd_net_),
            .in3(N__32301),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__47309),
            .ce(N__32404),
            .sr(N__46925));
    defparam \current_shift_inst.timer_s1.counter_17_LC_12_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_12_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_12_21_1  (
            .in0(N__33342),
            .in1(N__32290),
            .in2(_gnd_net_),
            .in3(N__32274),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__47309),
            .ce(N__32404),
            .sr(N__46925));
    defparam \current_shift_inst.timer_s1.counter_18_LC_12_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_12_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_12_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_12_21_2  (
            .in0(N__33312),
            .in1(N__32258),
            .in2(_gnd_net_),
            .in3(N__32244),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__47309),
            .ce(N__32404),
            .sr(N__46925));
    defparam \current_shift_inst.timer_s1.counter_19_LC_12_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_12_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_12_21_3  (
            .in0(N__33343),
            .in1(N__32228),
            .in2(_gnd_net_),
            .in3(N__32214),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__47309),
            .ce(N__32404),
            .sr(N__46925));
    defparam \current_shift_inst.timer_s1.counter_20_LC_12_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_12_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_12_21_4  (
            .in0(N__33313),
            .in1(N__32204),
            .in2(_gnd_net_),
            .in3(N__32190),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__47309),
            .ce(N__32404),
            .sr(N__46925));
    defparam \current_shift_inst.timer_s1.counter_21_LC_12_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_12_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_12_21_5  (
            .in0(N__33344),
            .in1(N__32185),
            .in2(_gnd_net_),
            .in3(N__32169),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__47309),
            .ce(N__32404),
            .sr(N__46925));
    defparam \current_shift_inst.timer_s1.counter_22_LC_12_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_12_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_12_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_12_21_6  (
            .in0(N__33314),
            .in1(N__32158),
            .in2(_gnd_net_),
            .in3(N__32142),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__47309),
            .ce(N__32404),
            .sr(N__46925));
    defparam \current_shift_inst.timer_s1.counter_23_LC_12_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_12_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_12_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_12_21_7  (
            .in0(N__33345),
            .in1(N__32579),
            .in2(_gnd_net_),
            .in3(N__32565),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__47309),
            .ce(N__32404),
            .sr(N__46925));
    defparam \current_shift_inst.timer_s1.counter_24_LC_12_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_12_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_12_22_0  (
            .in0(N__33336),
            .in1(N__32554),
            .in2(_gnd_net_),
            .in3(N__32538),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__47308),
            .ce(N__32412),
            .sr(N__46930));
    defparam \current_shift_inst.timer_s1.counter_25_LC_12_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_12_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_12_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_12_22_1  (
            .in0(N__33340),
            .in1(N__32524),
            .in2(_gnd_net_),
            .in3(N__32508),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__47308),
            .ce(N__32412),
            .sr(N__46930));
    defparam \current_shift_inst.timer_s1.counter_26_LC_12_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_12_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_12_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_12_22_2  (
            .in0(N__33337),
            .in1(N__32492),
            .in2(_gnd_net_),
            .in3(N__32478),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__47308),
            .ce(N__32412),
            .sr(N__46930));
    defparam \current_shift_inst.timer_s1.counter_27_LC_12_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_12_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_12_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_12_22_3  (
            .in0(N__33341),
            .in1(N__32473),
            .in2(_gnd_net_),
            .in3(N__32457),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__47308),
            .ce(N__32412),
            .sr(N__46930));
    defparam \current_shift_inst.timer_s1.counter_28_LC_12_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_12_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_12_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_12_22_4  (
            .in0(N__33338),
            .in1(N__32450),
            .in2(_gnd_net_),
            .in3(N__32436),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__47308),
            .ce(N__32412),
            .sr(N__46930));
    defparam \current_shift_inst.timer_s1.counter_29_LC_12_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_12_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_12_22_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_12_22_5  (
            .in0(N__32426),
            .in1(N__33339),
            .in2(_gnd_net_),
            .in3(N__32433),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47308),
            .ce(N__32412),
            .sr(N__46930));
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_12_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_12_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIC90O_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__33666),
            .in2(_gnd_net_),
            .in3(N__33744),
            .lcout(\current_shift_inst.timer_phase.N_188_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_7.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_7.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32640),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_13_4_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_13_4_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_13_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_13_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32616),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47427),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_13_5_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_13_5_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_13_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_13_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32598),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47420),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_6_0 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_6_0  (
            .in0(N__32745),
            .in1(N__36229),
            .in2(N__34017),
            .in3(N__32867),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(N__46813));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_13_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_13_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_13_6_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_13_6_1  (
            .in0(N__32864),
            .in1(N__32749),
            .in2(N__36245),
            .in3(N__33993),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(N__46813));
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_13_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_13_6_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_31_LC_13_6_2  (
            .in0(N__41879),
            .in1(N__40798),
            .in2(N__37841),
            .in3(N__39041),
            .lcout(measured_delay_hc_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(N__46813));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_6_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_6_3  (
            .in0(N__32861),
            .in1(N__32746),
            .in2(N__36242),
            .in3(N__33792),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(N__46813));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_6_4 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_6_4  (
            .in0(N__32744),
            .in1(N__36228),
            .in2(N__33756),
            .in3(N__32866),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(N__46813));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_6_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_6_5  (
            .in0(N__32862),
            .in1(N__32747),
            .in2(N__36243),
            .in3(N__34059),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(N__46813));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_13_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_13_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_13_6_6 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_13_6_6  (
            .in0(N__32743),
            .in1(N__36227),
            .in2(N__34128),
            .in3(N__32865),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(N__46813));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_6_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_6_7  (
            .in0(N__32863),
            .in1(N__32748),
            .in2(N__36244),
            .in3(N__34038),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(N__46813));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_7_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_7_0  (
            .in0(N__32736),
            .in1(N__32871),
            .in2(N__36234),
            .in3(N__34218),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47404),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_13_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_13_7_1 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_13_7_1  (
            .in0(N__32868),
            .in1(N__36197),
            .in2(N__33921),
            .in3(N__32740),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47404),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_7_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_7_2  (
            .in0(N__32737),
            .in1(N__32872),
            .in2(N__36235),
            .in3(N__34197),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47404),
            .ce(),
            .sr(N__46818));
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_13_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_13_7_3 .LUT_INIT=16'b1101100011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_6_LC_13_7_3  (
            .in0(N__40808),
            .in1(N__41259),
            .in2(N__36956),
            .in3(N__40916),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47404),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_13_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_13_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_13_7_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_13_7_4  (
            .in0(N__32739),
            .in1(N__32874),
            .in2(N__36237),
            .in3(N__33942),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47404),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_13_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_13_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_13_7_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_13_7_5  (
            .in0(N__32869),
            .in1(N__36198),
            .in2(N__34242),
            .in3(N__32741),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47404),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_13_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_13_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_13_7_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_13_7_6  (
            .in0(N__32738),
            .in1(N__32873),
            .in2(N__36236),
            .in3(N__34176),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47404),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_13_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_13_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_13_7_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_13_7_7  (
            .in0(N__32870),
            .in1(N__36199),
            .in2(N__34155),
            .in3(N__32742),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47404),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_13_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_13_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_13_8_0 .LUT_INIT=16'b1100100010001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_13_8_0  (
            .in0(N__32730),
            .in1(N__34083),
            .in2(N__36239),
            .in3(N__32860),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47395),
            .ce(),
            .sr(N__46822));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_13_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_13_8_1 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_13_8_1  (
            .in0(N__32856),
            .in1(N__36200),
            .in2(N__32761),
            .in3(N__34332),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47395),
            .ce(),
            .sr(N__46822));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_8_3 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_8_3  (
            .in0(N__32857),
            .in1(N__36201),
            .in2(N__32762),
            .in3(N__32901),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47395),
            .ce(),
            .sr(N__46822));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_13_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_13_8_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_13_8_4  (
            .in0(N__32729),
            .in1(N__32859),
            .in2(N__36238),
            .in3(N__34104),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47395),
            .ce(),
            .sr(N__46822));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_13_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_13_8_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_13_8_5  (
            .in0(N__32858),
            .in1(N__36202),
            .in2(N__32763),
            .in3(N__33969),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47395),
            .ce(),
            .sr(N__46822));
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_13_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_13_8_6 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_25_LC_13_8_6  (
            .in0(N__41637),
            .in1(N__40822),
            .in2(N__32894),
            .in3(N__40622),
            .lcout(measured_delay_hc_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47395),
            .ce(),
            .sr(N__46822));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_9_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_9_0  (
            .in0(N__32855),
            .in1(N__32731),
            .in2(N__36240),
            .in3(N__34581),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47385),
            .ce(N__34781),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__34626),
            .in2(_gnd_net_),
            .in3(N__34579),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_13_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_13_9_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_13_9_3  (
            .in0(N__34580),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34627),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_9_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_9_4  (
            .in0(N__47686),
            .in1(N__47514),
            .in2(N__47940),
            .in3(N__45968),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47385),
            .ce(N__34781),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_9_5 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_9_5  (
            .in0(N__45969),
            .in1(N__47932),
            .in2(N__47535),
            .in3(N__47687),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47385),
            .ce(N__34781),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_9_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_9_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_9_6  (
            .in0(N__44819),
            .in1(N__44622),
            .in2(N__42231),
            .in3(N__44696),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47385),
            .ce(N__34781),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_9_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_9_7 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_9_7  (
            .in0(N__44621),
            .in1(N__42226),
            .in2(N__44729),
            .in3(N__44820),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47385),
            .ce(N__34781),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_13_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_13_10_0 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_26_LC_13_10_0  (
            .in0(N__41961),
            .in1(N__40821),
            .in2(N__32967),
            .in3(N__40639),
            .lcout(measured_delay_hc_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47378),
            .ce(),
            .sr(N__46833));
    defparam \phase_controller_inst1.state_3_LC_13_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_13_10_2 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \phase_controller_inst1.state_3_LC_13_10_2  (
            .in0(N__34553),
            .in1(N__34656),
            .in2(N__34522),
            .in3(N__42029),
            .lcout(\phase_controller_inst1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47378),
            .ce(),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_13_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_13_10_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_13_10_3  (
            .in0(N__40640),
            .in1(N__40823),
            .in2(N__37233),
            .in3(N__41220),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47378),
            .ce(),
            .sr(N__46833));
    defparam \phase_controller_inst1.state_4_LC_13_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_13_10_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_13_10_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__35037),
            .in2(_gnd_net_),
            .in3(N__42055),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47378),
            .ce(),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_13_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_13_10_6 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_24_LC_13_10_6  (
            .in0(N__32948),
            .in1(N__40820),
            .in2(N__41894),
            .in3(N__39015),
            .lcout(measured_delay_hc_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47378),
            .ce(),
            .sr(N__46833));
    defparam \phase_controller_inst1.S1_LC_13_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34514),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47373),
            .ce(),
            .sr(N__46841));
    defparam \phase_controller_inst1.state_0_LC_13_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_13_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_13_11_4 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst1.state_0_LC_13_11_4  (
            .in0(N__42009),
            .in1(N__34683),
            .in2(N__34730),
            .in3(N__33044),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47373),
            .ce(),
            .sr(N__46841));
    defparam \current_shift_inst.timer_s1.running_LC_13_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_11_6 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_11_6  (
            .in0(N__33154),
            .in1(N__33369),
            .in2(_gnd_net_),
            .in3(N__33116),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47373),
            .ce(),
            .sr(N__46841));
    defparam \delay_measurement_inst.start_timer_hc_LC_13_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_13_12_2 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_13_12_2  (
            .in0(N__33088),
            .in1(N__33072),
            .in2(_gnd_net_),
            .in3(N__34287),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47365),
            .ce(),
            .sr(N__46844));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_13_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_13_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__42007),
            .in2(_gnd_net_),
            .in3(N__33040),
            .lcout(\phase_controller_inst1.N_231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.T01_sbtinv_LC_13_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_sbtinv_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.T01_sbtinv_LC_13_13_0 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \phase_controller_inst1.T01_sbtinv_LC_13_13_0  (
            .in0(N__42008),
            .in1(N__34729),
            .in2(N__34526),
            .in3(N__33045),
            .lcout(\phase_controller_inst1.N_221_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync1_LC_13_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync1_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync1_LC_13_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S3_sync1_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33000),
            .lcout(\current_shift_inst.S3_syncZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47357),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_13_13_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_13_13_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_13_13_5  (
            .in0(N__42115),
            .in1(N__44821),
            .in2(_gnd_net_),
            .in3(N__44707),
            .lcout(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_13_13_6 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_13_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_0_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__34876),
            .in2(_gnd_net_),
            .in3(N__34857),
            .lcout(\phase_controller_slave.N_214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync0_LC_13_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync0_LC_13_13_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync0_LC_13_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.S3_sync0_LC_13_13_7  (
            .in0(N__34819),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.S3_syncZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47357),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32994),
            .lcout(\current_shift_inst.un4_control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32973),
            .lcout(\current_shift_inst.un4_control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33408),
            .lcout(\current_shift_inst.un4_control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33390),
            .lcout(\current_shift_inst.un4_control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33372),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_14_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_14_6  (
            .in0(N__33213),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_14_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_14_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(N__45660),
            .in2(_gnd_net_),
            .in3(N__45363),
            .lcout(\phase_controller_slave.stoper_tr.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_13_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_13_15_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_13_15_1  (
            .in0(N__47900),
            .in1(N__47725),
            .in2(_gnd_net_),
            .in3(N__47542),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33192),
            .lcout(\current_shift_inst.un4_control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__33174),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33510),
            .lcout(\current_shift_inst.un4_control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33492),
            .lcout(\current_shift_inst.un4_control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_13_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_13_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_13_16_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_13_16_1  (
            .in0(N__42680),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43156),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47334),
            .ce(N__43046),
            .sr(N__46882));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_13_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_13_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_13_16_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_13_16_2  (
            .in0(N__43157),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42647),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47334),
            .ce(N__43046),
            .sr(N__46882));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_13_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_13_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_13_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__43158),
            .in2(_gnd_net_),
            .in3(N__42611),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47334),
            .ce(N__43046),
            .sr(N__46882));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33474),
            .lcout(\current_shift_inst.un4_control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33456),
            .lcout(\current_shift_inst.un4_control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33438),
            .lcout(\current_shift_inst.un4_control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_13_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_13_17_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__46984),
            .in2(_gnd_net_),
            .in3(N__39602),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_17_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_17_1  (
            .in0(N__35627),
            .in1(N__33525),
            .in2(N__38075),
            .in3(N__33584),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_13_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_13_17_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_13_17_2  (
            .in0(N__39669),
            .in1(N__33900),
            .in2(N__33540),
            .in3(N__35237),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_321_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_13_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_13_17_3 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_13_17_3  (
            .in0(N__35238),
            .in1(N__36433),
            .in2(N__33537),
            .in3(N__33531),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_13_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_13_17_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_13_17_4  (
            .in0(N__33585),
            .in1(N__35942),
            .in2(N__33519),
            .in3(N__35970),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_13_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_13_17_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_13_17_5  (
            .in0(N__33555),
            .in1(N__35750),
            .in2(N__33534),
            .in3(N__35820),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_13_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_13_17_7 .LUT_INIT=16'b0000000011110100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_13_17_7  (
            .in0(N__33901),
            .in1(N__39670),
            .in2(N__35295),
            .in3(N__36434),
            .lcout(\delay_measurement_inst.N_284_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_18_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_18_0  (
            .in0(N__35741),
            .in1(N__35639),
            .in2(N__35459),
            .in3(N__35817),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_18_1  (
            .in0(N__38289),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47323),
            .ce(N__36365),
            .sr(N__46902));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38262),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47323),
            .ce(N__36365),
            .sr(N__46902));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_13_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_13_18_3 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_13_18_3  (
            .in0(N__35906),
            .in1(N__35452),
            .in2(N__35883),
            .in3(N__35626),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_13_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_13_18_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__35837),
            .in2(_gnd_net_),
            .in3(N__35435),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_320_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_13_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_13_18_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_13_18_6  (
            .in0(N__35966),
            .in1(N__35882),
            .in2(N__35943),
            .in3(N__35907),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_13_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_13_19_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_13_19_1 .LUT_INIT=16'b0011000000110001;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_13_19_1  (
            .in0(N__33572),
            .in1(N__33870),
            .in2(N__35749),
            .in3(N__36439),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47319),
            .ce(N__35508),
            .sr(N__46909));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_13_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_13_19_2 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_13_19_2  (
            .in0(N__33554),
            .in1(N__33902),
            .in2(_gnd_net_),
            .in3(N__35290),
            .lcout(\delay_measurement_inst.N_305_1 ),
            .ltout(\delay_measurement_inst.N_305_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_13_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_13_19_3 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__36437),
            .in2(N__33576),
            .in3(N__35703),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47319),
            .ce(N__35508),
            .sr(N__46909));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_13_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_13_19_4 .LUT_INIT=16'b1010100010101000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_13_19_4  (
            .in0(N__35688),
            .in1(N__33567),
            .in2(N__36454),
            .in3(_gnd_net_),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47319),
            .ce(N__35508),
            .sr(N__46909));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_13_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_13_19_5 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__36438),
            .in2(N__33573),
            .in3(N__35667),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47319),
            .ce(N__35508),
            .sr(N__46909));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_13_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_13_19_6 .LUT_INIT=16'b1010100010101000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_13_19_6  (
            .in0(N__36003),
            .in1(N__33571),
            .in2(N__36455),
            .in3(_gnd_net_),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47319),
            .ce(N__35508),
            .sr(N__46909));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_13_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_13_20_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_13_20_0 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_13_20_0  (
            .in0(N__36432),
            .in1(N__35878),
            .in2(_gnd_net_),
            .in3(N__35288),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47316),
            .ce(N__35507),
            .sr(N__46915));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_13_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_13_20_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__39643),
            .in2(_gnd_net_),
            .in3(N__38056),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_13_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_13_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_13_21_3  (
            .in0(N__33591),
            .in1(N__33597),
            .in2(N__35856),
            .in3(N__33879),
            .lcout(\delay_measurement_inst.N_358 ),
            .ltout(\delay_measurement_inst.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_13_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_13_21_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_13_21_4 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__36430),
            .in2(N__33747),
            .in3(N__35965),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47313),
            .ce(N__35509),
            .sr(N__46922));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_13_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_13_21_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_13_21_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_13_21_5  (
            .in0(N__36429),
            .in1(N__35932),
            .in2(_gnd_net_),
            .in3(N__35287),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47313),
            .ce(N__35509),
            .sr(N__46922));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_13_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_13_21_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_13_21_6  (
            .in0(N__35286),
            .in1(N__36431),
            .in2(_gnd_net_),
            .in3(N__35900),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47313),
            .ce(N__35509),
            .sr(N__46922));
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_13_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_13_22_0 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIL91O_LC_13_22_0  (
            .in0(N__33742),
            .in1(N__33701),
            .in2(_gnd_net_),
            .in3(N__33675),
            .lcout(\current_shift_inst.timer_phase.N_192_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_13_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_13_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_13_22_2  (
            .in0(N__36033),
            .in1(N__36042),
            .in2(N__36024),
            .in3(N__36051),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__35343),
            .in2(_gnd_net_),
            .in3(N__39981),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_337_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_13_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_13_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_13_22_4  (
            .in0(N__36072),
            .in1(N__36081),
            .in2(N__36063),
            .in3(N__35844),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_13_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_13_22_5 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_13_22_5  (
            .in0(N__35745),
            .in1(N__38062),
            .in2(_gnd_net_),
            .in3(N__35591),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_13_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_13_22_6 .LUT_INIT=16'b0000000011011100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_13_22_6  (
            .in0(N__39653),
            .in1(N__33909),
            .in2(N__33882),
            .in3(N__35285),
            .lcout(\delay_measurement_inst.N_324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_13_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_13_23_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__36468),
            .in2(_gnd_net_),
            .in3(N__36012),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_13_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_13_23_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_13_23_5  (
            .in0(N__35592),
            .in1(N__39671),
            .in2(N__35751),
            .in3(N__35294),
            .lcout(\delay_measurement_inst.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_28_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_28_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_28_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_28_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34734),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(),
            .sr(N__46945));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_1  (
            .in0(_gnd_net_),
            .in1(N__40954),
            .in2(_gnd_net_),
            .in3(N__43000),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_335_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_4_2  (
            .in0(_gnd_net_),
            .in1(N__34527),
            .in2(_gnd_net_),
            .in3(N__34546),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_14_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_14_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(N__33840),
            .in2(N__33828),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_14_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_14_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__33804),
            .in2(_gnd_net_),
            .in3(N__33786),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_14_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_14_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__33783),
            .in2(N__33771),
            .in3(N__34074),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_14_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_14_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(N__34071),
            .in2(_gnd_net_),
            .in3(N__34053),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_14_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_14_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(N__34050),
            .in2(_gnd_net_),
            .in3(N__34032),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_14_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_14_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(N__34029),
            .in2(_gnd_net_),
            .in3(N__34008),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_14_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_14_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(N__34005),
            .in2(_gnd_net_),
            .in3(N__33987),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_14_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_14_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__33984),
            .in2(_gnd_net_),
            .in3(N__33957),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_14_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_14_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(N__33954),
            .in2(_gnd_net_),
            .in3(N__33936),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_14_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_14_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__33933),
            .in2(_gnd_net_),
            .in3(N__33912),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_14_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_14_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__34254),
            .in2(_gnd_net_),
            .in3(N__34233),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_14_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_14_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__34230),
            .in2(_gnd_net_),
            .in3(N__34212),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_14_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_14_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__34209),
            .in2(_gnd_net_),
            .in3(N__34191),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_14_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_14_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__34188),
            .in2(_gnd_net_),
            .in3(N__34170),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_14_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_14_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(N__34167),
            .in2(_gnd_net_),
            .in3(N__34146),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_14_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_14_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__34142),
            .in2(_gnd_net_),
            .in3(N__34119),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_14_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_14_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__34116),
            .in2(_gnd_net_),
            .in3(N__34098),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_14_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_14_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__34095),
            .in2(_gnd_net_),
            .in3(N__34077),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_14_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_14_7_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__34347),
            .in2(_gnd_net_),
            .in3(N__34335),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_7_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__36857),
            .in2(_gnd_net_),
            .in3(N__40878),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_a3_LC_14_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_a3_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_a3_LC_14_7_4 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m3_0_a3_LC_14_7_4  (
            .in0(N__37037),
            .in1(N__36938),
            .in2(N__34326),
            .in3(N__34311),
            .lcout(\phase_controller_inst1.stoper_hc.un1_N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_7_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_7_5  (
            .in0(N__39006),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41824),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_14_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_14_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_14_7_6  (
            .in0(N__36826),
            .in1(N__36899),
            .in2(N__37739),
            .in3(N__36978),
            .lcout(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__34473),
            .in2(_gnd_net_),
            .in3(N__34449),
            .lcout(\phase_controller_inst1.N_228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_14_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_14_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_14_8_1  (
            .in0(N__36590),
            .in1(N__36630),
            .in2(N__37550),
            .in3(N__36683),
            .lcout(\phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_14_8_5.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_14_8_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_14_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_14_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41004),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47405),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_8_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__41853),
            .in2(_gnd_net_),
            .in3(N__39005),
            .lcout(\delay_measurement_inst.delay_hc_reg3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_1_LC_14_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_14_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_14_9_0 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst1.state_1_LC_14_9_0  (
            .in0(N__34681),
            .in1(N__34451),
            .in2(N__34725),
            .in3(N__34476),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47396),
            .ce(),
            .sr(N__46823));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_14_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_14_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_14_9_1 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_14_9_1  (
            .in0(N__34475),
            .in1(N__34638),
            .in2(N__34605),
            .in3(N__34590),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47396),
            .ce(),
            .sr(N__46823));
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_14_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_14_9_2 .LUT_INIT=16'b1111111010111010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_14_LC_14_9_2  (
            .in0(N__40618),
            .in1(N__40811),
            .in2(N__36750),
            .in3(N__41496),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47396),
            .ce(),
            .sr(N__46823));
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_14_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_14_9_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_13_LC_14_9_3  (
            .in0(N__40809),
            .in1(N__41523),
            .in2(N__37560),
            .in3(N__40617),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47396),
            .ce(),
            .sr(N__46823));
    defparam \delay_measurement_inst.prev_tr_sig_LC_14_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_tr_sig_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_tr_sig_LC_14_9_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.prev_tr_sig_LC_14_9_4  (
            .in0(N__36303),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.prev_tr_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47396),
            .ce(),
            .sr(N__46823));
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_14_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_14_9_5 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_18_LC_14_9_5  (
            .in0(N__40810),
            .in1(N__41730),
            .in2(N__34426),
            .in3(N__40619),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47396),
            .ce(),
            .sr(N__46823));
    defparam \phase_controller_inst1.state_2_LC_14_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_14_9_6 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_14_9_6  (
            .in0(N__34554),
            .in1(N__34450),
            .in2(N__34521),
            .in3(N__34474),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47396),
            .ce(),
            .sr(N__46823));
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_2 .LUT_INIT=16'b1111000000010000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_2  (
            .in0(N__34383),
            .in1(N__37865),
            .in2(N__37439),
            .in3(N__34415),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(N__37091),
            .sr(N__46828));
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_10_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_12_LC_14_10_6  (
            .in0(N__36607),
            .in1(N__37186),
            .in2(N__37440),
            .in3(N__37495),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(N__37091),
            .sr(N__46828));
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_7 .LUT_INIT=16'b1000100010001100;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_7  (
            .in0(N__36500),
            .in1(N__37429),
            .in2(N__37883),
            .in3(N__34382),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(N__37091),
            .sr(N__46828));
    defparam reset_ibuf_gb_io_RNI79U7_LC_14_11_0.C_ON=1'b0;
    defparam reset_ibuf_gb_io_RNI79U7_LC_14_11_0.SEQ_MODE=4'b0000;
    defparam reset_ibuf_gb_io_RNI79U7_LC_14_11_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 reset_ibuf_gb_io_RNI79U7_LC_14_11_0 (
            .in0(N__46977),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(red_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__34718),
            .in2(_gnd_net_),
            .in3(N__34682),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_11_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_11_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_11_6  (
            .in0(N__42130),
            .in1(N__44822),
            .in2(_gnd_net_),
            .in3(N__44708),
            .lcout(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_14_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_14_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__35054),
            .in2(_gnd_net_),
            .in3(N__42054),
            .lcout(\phase_controller_inst1.N_232 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_14_12_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_14_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_14_12_6 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_9_LC_14_12_6  (
            .in0(N__37411),
            .in1(N__37042),
            .in2(_gnd_net_),
            .in3(N__37690),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__37099),
            .sr(N__46842));
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_14_12_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_14_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_14_12_7 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_19_LC_14_12_7  (
            .in0(N__37691),
            .in1(N__37881),
            .in2(_gnd_net_),
            .in3(N__36558),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__37099),
            .sr(N__46842));
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_14_13_0 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_14_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_1_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__35161),
            .in2(_gnd_net_),
            .in3(N__35197),
            .lcout(\phase_controller_slave.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_2_LC_14_13_3 .C_ON=1'b0;
    defparam \phase_controller_slave.state_2_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_2_LC_14_13_3 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_slave.state_2_LC_14_13_3  (
            .in0(N__35198),
            .in1(N__34877),
            .in2(N__35166),
            .in3(N__34858),
            .lcout(\phase_controller_slave.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47366),
            .ce(),
            .sr(N__46845));
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_14_13_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_14_13_5 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_LC_14_13_5  (
            .in0(N__34859),
            .in1(N__44649),
            .in2(N__34650),
            .in3(N__44620),
            .lcout(\phase_controller_slave.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47366),
            .ce(),
            .sr(N__46845));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_13_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_13_6 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_13_6  (
            .in0(N__44873),
            .in1(N__42129),
            .in2(N__44772),
            .in3(N__44406),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47366),
            .ce(),
            .sr(N__46845));
    defparam \phase_controller_slave.start_timer_hc_LC_14_14_0 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_LC_14_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_hc_LC_14_14_0 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_slave.start_timer_hc_LC_14_14_0  (
            .in0(N__34942),
            .in1(N__34914),
            .in2(N__42192),
            .in3(N__34908),
            .lcout(\phase_controller_slave.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47358),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_slave.S2_LC_14_14_2 .C_ON=1'b0;
    defparam \phase_controller_slave.S2_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S2_LC_14_14_2 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \phase_controller_slave.S2_LC_14_14_2  (
            .in0(N__34974),
            .in1(N__35157),
            .in2(N__34895),
            .in3(N__35406),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47358),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_slave.state_1_LC_14_14_3 .C_ON=1'b0;
    defparam \phase_controller_slave.state_1_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_1_LC_14_14_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_slave.state_1_LC_14_14_3  (
            .in0(N__35385),
            .in1(N__34878),
            .in2(N__35412),
            .in3(N__34860),
            .lcout(\phase_controller_slave.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47358),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_slave.S1_LC_14_14_4 .C_ON=1'b0;
    defparam \phase_controller_slave.S1_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S1_LC_14_14_4 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \phase_controller_slave.S1_LC_14_14_4  (
            .in0(N__34973),
            .in1(_gnd_net_),
            .in2(N__34823),
            .in3(N__35156),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47358),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_slave.state_4_LC_14_14_5 .C_ON=1'b0;
    defparam \phase_controller_slave.state_4_LC_14_14_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.state_4_LC_14_14_5 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_slave.state_4_LC_14_14_5  (
            .in0(N__35055),
            .in1(N__34972),
            .in2(_gnd_net_),
            .in3(N__34941),
            .lcout(\phase_controller_slave.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47358),
            .ce(),
            .sr(N__46853));
    defparam \delay_measurement_inst.start_timer_tr_LC_14_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_14_14_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_14_14_6 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_14_14_6  (
            .in0(N__36291),
            .in1(N__35132),
            .in2(_gnd_net_),
            .in3(N__35101),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47358),
            .ce(),
            .sr(N__46853));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_14_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_14_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_14_14_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_14_14_7  (
            .in0(N__35339),
            .in1(N__35312),
            .in2(_gnd_net_),
            .in3(N__39976),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47358),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_14_15_0 .C_ON=1'b0;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_14_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.state_RNIVDE2_0_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__35218),
            .in2(_gnd_net_),
            .in3(N__35207),
            .lcout(\phase_controller_slave.N_211 ),
            .ltout(\phase_controller_slave.N_211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_tr_LC_14_15_1 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_tr_LC_14_15_1 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_slave.start_timer_tr_LC_14_15_1  (
            .in0(N__45533),
            .in1(N__35352),
            .in2(N__34800),
            .in3(N__34943),
            .lcout(\phase_controller_slave.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(),
            .sr(N__46862));
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_14_15_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_14_15_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_14_15_2  (
            .in0(N__45495),
            .in1(N__45730),
            .in2(_gnd_net_),
            .in3(N__45411),
            .lcout(),
            .ltout(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_14_15_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_14_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_14_15_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_LC_14_15_3  (
            .in0(N__35222),
            .in1(N__39528),
            .in2(N__35226),
            .in3(N__41091),
            .lcout(\phase_controller_slave.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(),
            .sr(N__46862));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_14_15_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_14_15_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_16_LC_14_15_4  (
            .in0(N__45723),
            .in1(N__45412),
            .in2(N__45534),
            .in3(N__37980),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(),
            .sr(N__46862));
    defparam \phase_controller_slave.state_0_LC_14_15_5 .C_ON=1'b0;
    defparam \phase_controller_slave.state_0_LC_14_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_0_LC_14_15_5 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_slave.state_0_LC_14_15_5  (
            .in0(N__35208),
            .in1(N__35410),
            .in2(N__35223),
            .in3(N__35384),
            .lcout(\phase_controller_slave.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(),
            .sr(N__46862));
    defparam \phase_controller_slave.state_3_LC_14_15_6 .C_ON=1'b0;
    defparam \phase_controller_slave.state_3_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_3_LC_14_15_6 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \phase_controller_slave.state_3_LC_14_15_6  (
            .in0(N__34920),
            .in1(N__35199),
            .in2(N__35165),
            .in3(N__35172),
            .lcout(\phase_controller_slave.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(),
            .sr(N__46862));
    defparam \delay_measurement_inst.stop_timer_tr_LC_14_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_14_16_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_14_16_6  (
            .in0(N__36301),
            .in1(N__35133),
            .in2(N__46989),
            .in3(N__35102),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47342),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_RNO_0_3_LC_14_16_7 .C_ON=1'b0;
    defparam \phase_controller_slave.state_RNO_0_3_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_RNO_0_3_LC_14_16_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.state_RNO_0_3_LC_14_16_7  (
            .in0(N__35065),
            .in1(N__34971),
            .in2(_gnd_net_),
            .in3(N__34944),
            .lcout(\phase_controller_slave.N_213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_14_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_14_17_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_14_17_0  (
            .in0(N__43259),
            .in1(N__46214),
            .in2(_gnd_net_),
            .in3(N__46174),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_14_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_14_17_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__43328),
            .in2(N__35415),
            .in3(N__42739),
            .lcout(\phase_controller_inst1.stoper_tr.N_20_li ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_14_17_2 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_14_17_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_tr_RNO_0_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__35411),
            .in2(_gnd_net_),
            .in3(N__35383),
            .lcout(\phase_controller_slave.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_17_3 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_17_3  (
            .in0(N__35332),
            .in1(N__35313),
            .in2(_gnd_net_),
            .in3(N__39972),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_338_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_14_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_14_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_14_17_4  (
            .in0(N__42646),
            .in1(N__42679),
            .in2(N__42612),
            .in3(N__43105),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_14_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_14_17_5 .LUT_INIT=16'b0000000001110101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_14_17_5  (
            .in0(N__42893),
            .in1(N__46255),
            .in2(N__35298),
            .in3(N__43258),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_14_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_14_18_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_5_LC_14_18_0  (
            .in0(N__35607),
            .in1(N__36448),
            .in2(N__35563),
            .in3(N__35838),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47328),
            .ce(N__35510),
            .sr(N__46889));
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_14_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_14_18_1 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_14_18_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_3_LC_14_18_1  (
            .in0(N__36447),
            .in1(N__35610),
            .in2(N__35460),
            .in3(N__35557),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47328),
            .ce(N__35510),
            .sr(N__46889));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_14_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_14_18_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_14_18_2  (
            .in0(N__35790),
            .in1(N__35576),
            .in2(N__35772),
            .in3(N__35289),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_331 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_14_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_14_18_3 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__39665),
            .in2(N__35229),
            .in3(N__35818),
            .lcout(\delay_measurement_inst.N_333 ),
            .ltout(\delay_measurement_inst.N_333_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_14_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_14_18_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_4_LC_14_18_4  (
            .in0(N__35549),
            .in1(N__35436),
            .in2(N__35643),
            .in3(N__36452),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47328),
            .ce(N__35510),
            .sr(N__46889));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_14_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_14_18_5 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_14_18_5  (
            .in0(N__36446),
            .in1(N__35608),
            .in2(N__35565),
            .in3(N__35819),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47328),
            .ce(N__35510),
            .sr(N__46889));
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_14_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_14_18_6 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_14_18_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_1_LC_14_18_6  (
            .in0(N__35609),
            .in1(N__35640),
            .in2(N__35564),
            .in3(N__36453),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47328),
            .ce(N__35510),
            .sr(N__46889));
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_14_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_14_18_7 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_2_LC_14_18_7  (
            .in0(N__35628),
            .in1(N__35550),
            .in2(N__36456),
            .in3(N__35606),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47328),
            .ce(N__35510),
            .sr(N__46889));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_19_0  (
            .in0(N__35663),
            .in1(N__35687),
            .in2(N__36002),
            .in3(N__35702),
            .lcout(\delay_measurement_inst.N_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_7_LC_14_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_7_LC_14_19_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_7_LC_14_19_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_7_LC_14_19_2  (
            .in0(N__36435),
            .in1(N__35561),
            .in2(_gnd_net_),
            .in3(N__35789),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47324),
            .ce(N__35511),
            .sr(N__46903));
    defparam \delay_measurement_inst.delay_tr_reg_esr_8_LC_14_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_8_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_8_LC_14_19_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_8_LC_14_19_4  (
            .in0(N__36436),
            .in1(N__35562),
            .in2(_gnd_net_),
            .in3(N__35768),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47324),
            .ce(N__35511),
            .sr(N__46903));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_14_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_14_19_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_14_19_5  (
            .in0(N__39574),
            .in1(N__42493),
            .in2(_gnd_net_),
            .in3(N__42844),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_20_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__38282),
            .in2(N__38235),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47320),
            .ce(N__36366),
            .sr(N__46910));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__38255),
            .in2(N__38211),
            .in3(N__35418),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47320),
            .ce(N__36366),
            .sr(N__46910));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__38234),
            .in2(N__38187),
            .in3(N__35823),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47320),
            .ce(N__36366),
            .sr(N__46910));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__38210),
            .in2(N__38163),
            .in3(N__35793),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47320),
            .ce(N__36366),
            .sr(N__46910));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__38186),
            .in2(N__38139),
            .in3(N__35775),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47320),
            .ce(N__36366),
            .sr(N__46910));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__38162),
            .in2(N__38505),
            .in3(N__35754),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47320),
            .ce(N__36366),
            .sr(N__46910));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__38138),
            .in2(N__38481),
            .in3(N__35706),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47320),
            .ce(N__36366),
            .sr(N__46910));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__38504),
            .in2(N__38457),
            .in3(N__35691),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47320),
            .ce(N__36366),
            .sr(N__46910));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__38480),
            .in2(N__38433),
            .in3(N__35670),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47317),
            .ce(N__36347),
            .sr(N__46916));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__38456),
            .in2(N__38409),
            .in3(N__35646),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47317),
            .ce(N__36347),
            .sr(N__46916));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__38432),
            .in2(N__38385),
            .in3(N__35979),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47317),
            .ce(N__36347),
            .sr(N__46916));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__38408),
            .in2(N__38361),
            .in3(N__35976),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47317),
            .ce(N__36347),
            .sr(N__46916));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__38384),
            .in2(N__38337),
            .in3(N__35973),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47317),
            .ce(N__36347),
            .sr(N__46916));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__38360),
            .in2(N__38313),
            .in3(N__35946),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47317),
            .ce(N__36347),
            .sr(N__46916));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__38336),
            .in2(N__38697),
            .in3(N__35910),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47317),
            .ce(N__36347),
            .sr(N__46916));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__38312),
            .in2(N__38673),
            .in3(N__35886),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47317),
            .ce(N__36347),
            .sr(N__46916));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(N__38696),
            .in2(N__38649),
            .in3(N__35859),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47314),
            .ce(N__36355),
            .sr(N__46923));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(N__38672),
            .in2(N__38625),
            .in3(N__35847),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47314),
            .ce(N__36355),
            .sr(N__46923));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(N__38648),
            .in2(N__38601),
            .in3(N__36084),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47314),
            .ce(N__36355),
            .sr(N__46923));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(N__38624),
            .in2(N__38577),
            .in3(N__36075),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47314),
            .ce(N__36355),
            .sr(N__46923));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__38600),
            .in2(N__38553),
            .in3(N__36066),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47314),
            .ce(N__36355),
            .sr(N__46923));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_22_5  (
            .in0(_gnd_net_),
            .in1(N__38576),
            .in2(N__38529),
            .in3(N__36054),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47314),
            .ce(N__36355),
            .sr(N__46923));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_22_6  (
            .in0(_gnd_net_),
            .in1(N__38552),
            .in2(N__38871),
            .in3(N__36045),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47314),
            .ce(N__36355),
            .sr(N__46923));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(N__38528),
            .in2(N__38847),
            .in3(N__36036),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47314),
            .ce(N__36355),
            .sr(N__46923));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__38870),
            .in2(N__38823),
            .in3(N__36027),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47311),
            .ce(N__36348),
            .sr(N__46926));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_23_1  (
            .in0(_gnd_net_),
            .in1(N__38846),
            .in2(N__38799),
            .in3(N__36015),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47311),
            .ce(N__36348),
            .sr(N__46926));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(N__38822),
            .in2(N__38775),
            .in3(N__36006),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47311),
            .ce(N__36348),
            .sr(N__46926));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(N__38798),
            .in2(N__38754),
            .in3(N__36462),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47311),
            .ce(N__36348),
            .sr(N__46926));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36459),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47311),
            .ce(N__36348),
            .sr(N__46926));
    defparam SB_DFF_inst_DELAY_TR1_LC_15_4_1.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_4_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_15_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36318),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47443),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR2_LC_15_4_2.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_4_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_15_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36309),
            .lcout(delay_tr_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47443),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_15_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_15_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_15_5_1 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_15_5_1  (
            .in0(N__36261),
            .in1(N__42072),
            .in2(N__36178),
            .in3(N__36255),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47436),
            .ce(),
            .sr(N__46804));
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_15_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_15_6_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_15_6_2 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_0_LC_15_6_2  (
            .in0(N__40784),
            .in1(N__36985),
            .in2(N__41899),
            .in3(N__39030),
            .lcout(measured_delay_hc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47428),
            .ce(),
            .sr(N__46807));
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_15_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_15_6_3 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_15_6_3 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_3_LC_15_6_3  (
            .in0(N__36867),
            .in1(N__40786),
            .in2(N__41346),
            .in3(N__40912),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47428),
            .ce(),
            .sr(N__46807));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6  (
            .in0(N__40989),
            .in1(N__40958),
            .in2(_gnd_net_),
            .in3(N__42999),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47428),
            .ce(),
            .sr(N__46807));
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_15_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_15_6_7 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_15_6_7 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_1_LC_15_6_7  (
            .in0(N__36909),
            .in1(N__40785),
            .in2(N__41388),
            .in3(N__40911),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47428),
            .ce(),
            .sr(N__46807));
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_15_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_15_7_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_5_LC_15_7_1  (
            .in0(N__40743),
            .in1(N__41289),
            .in2(N__37747),
            .in3(N__40630),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47421),
            .ce(),
            .sr(N__46810));
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_15_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_15_7_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_11_LC_15_7_3  (
            .in0(N__40742),
            .in1(N__41583),
            .in2(N__36648),
            .in3(N__40628),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47421),
            .ce(),
            .sr(N__46810));
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_15_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_15_7_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_15_7_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_12_LC_15_7_4  (
            .in0(N__40629),
            .in1(N__40744),
            .in2(N__36608),
            .in3(N__41553),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47421),
            .ce(),
            .sr(N__46810));
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_15_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_15_8_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_15_8_4 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_19_LC_15_8_4  (
            .in0(N__40775),
            .in1(N__41709),
            .in2(N__36551),
            .in3(N__40620),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47414),
            .ce(),
            .sr(N__46814));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_15_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_15_8_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_15_8_7  (
            .in0(N__40621),
            .in1(N__40776),
            .in2(N__37932),
            .in3(N__41187),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47414),
            .ce(),
            .sr(N__46814));
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_15_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_15_9_1 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_4_LC_15_9_1  (
            .in0(N__36825),
            .in1(N__40777),
            .in2(N__41319),
            .in3(N__40626),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47406),
            .ce(),
            .sr(N__46819));
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_15_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_15_9_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_15_9_2 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_17_LC_15_9_2  (
            .in0(N__40625),
            .in1(N__36501),
            .in2(N__40819),
            .in3(N__41409),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47406),
            .ce(),
            .sr(N__46819));
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_15_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_15_9_5 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_10_LC_15_9_5  (
            .in0(N__36693),
            .in1(N__41613),
            .in2(N__40832),
            .in3(N__40623),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47406),
            .ce(),
            .sr(N__46819));
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_15_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_15_9_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_15_9_6 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_16_LC_15_9_6  (
            .in0(N__40624),
            .in1(N__36775),
            .in2(N__40818),
            .in3(N__41433),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47406),
            .ce(),
            .sr(N__46819));
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_15_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_15_9_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_15_9_7 .LUT_INIT=16'b1111111111001010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_9_LC_15_9_7  (
            .in0(N__37036),
            .in1(N__41154),
            .in2(N__40833),
            .in3(N__40627),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47406),
            .ce(),
            .sr(N__46819));
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_15_10_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_15_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_15_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_0_LC_15_10_0  (
            .in0(N__37187),
            .in1(N__37508),
            .in2(N__36993),
            .in3(N__37428),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47397),
            .ce(N__37106),
            .sr(N__46824));
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_10_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_10_1 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_10_1  (
            .in0(N__37421),
            .in1(N__36957),
            .in2(_gnd_net_),
            .in3(N__37645),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47397),
            .ce(N__37106),
            .sr(N__46824));
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_15_10_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_15_10_2 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_1_LC_15_10_2  (
            .in0(N__37647),
            .in1(N__37423),
            .in2(_gnd_net_),
            .in3(N__36914),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47397),
            .ce(N__37106),
            .sr(N__46824));
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_15_10_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_15_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_15_10_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_2_LC_15_10_3  (
            .in0(N__40885),
            .in1(_gnd_net_),
            .in2(N__37438),
            .in3(N__37648),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47397),
            .ce(N__37106),
            .sr(N__46824));
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_15_10_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_15_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_15_10_4 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_3_LC_15_10_4  (
            .in0(N__37649),
            .in1(N__37424),
            .in2(_gnd_net_),
            .in3(N__36876),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47397),
            .ce(N__37106),
            .sr(N__46824));
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_15_10_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_15_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_15_10_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_4_LC_15_10_5  (
            .in0(N__37882),
            .in1(N__36824),
            .in2(_gnd_net_),
            .in3(N__37650),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47397),
            .ce(N__37106),
            .sr(N__46824));
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_15_10_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_15_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_15_10_7 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_16_LC_15_10_7  (
            .in0(N__37422),
            .in1(N__36774),
            .in2(_gnd_net_),
            .in3(N__37646),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47397),
            .ce(N__37106),
            .sr(N__46824));
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_15_11_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_15_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_15_11_0 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_14_LC_15_11_0  (
            .in0(N__36749),
            .in1(_gnd_net_),
            .in2(N__37436),
            .in3(N__37681),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47387),
            .ce(N__37092),
            .sr(N__46829));
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_15_11_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_15_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_15_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_10_LC_15_11_2  (
            .in0(N__36697),
            .in1(N__37188),
            .in2(N__37437),
            .in3(N__37509),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47387),
            .ce(N__37092),
            .sr(N__46829));
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_15_11_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_15_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_15_11_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_8_LC_15_11_3  (
            .in0(N__37683),
            .in1(N__37887),
            .in2(_gnd_net_),
            .in3(N__37928),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47387),
            .ce(N__37092),
            .sr(N__46829));
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_15_11_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_15_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_15_11_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_5_LC_15_11_4  (
            .in0(N__37886),
            .in1(N__37743),
            .in2(_gnd_net_),
            .in3(N__37682),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47387),
            .ce(N__37092),
            .sr(N__46829));
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_15_11_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_15_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_15_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_13_LC_15_11_5  (
            .in0(N__37510),
            .in1(N__37416),
            .in2(N__37562),
            .in3(N__37190),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47387),
            .ce(N__37092),
            .sr(N__46829));
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_15_11_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_15_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_15_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_15_LC_15_11_6  (
            .in0(N__37412),
            .in1(N__37189),
            .in2(N__40562),
            .in3(N__37511),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47387),
            .ce(N__37092),
            .sr(N__46829));
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_15_11_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_15_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_15_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_7_LC_15_11_7  (
            .in0(N__37512),
            .in1(N__37417),
            .in2(N__37241),
            .in3(N__37191),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47387),
            .ce(N__37092),
            .sr(N__46829));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_0  (
            .in0(N__47721),
            .in1(N__47570),
            .in2(N__47939),
            .in3(N__45060),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47379),
            .ce(),
            .sr(N__46834));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_12_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_12_1  (
            .in0(N__47569),
            .in1(N__47926),
            .in2(N__47741),
            .in3(N__45021),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47379),
            .ce(),
            .sr(N__46834));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_12_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_12_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_12_3  (
            .in0(N__44891),
            .in1(N__44751),
            .in2(N__42230),
            .in3(N__39378),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47379),
            .ce(),
            .sr(N__46834));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_12_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_12_6 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_12_6  (
            .in0(N__44750),
            .in1(N__44892),
            .in2(N__44469),
            .in3(N__42217),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47379),
            .ce(),
            .sr(N__46834));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__39540),
            .in2(N__39801),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_15_13_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_15_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__39762),
            .in2(_gnd_net_),
            .in3(N__37965),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_15_13_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_15_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__39504),
            .in2(N__39738),
            .in3(N__37962),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_15_13_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_15_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__40296),
            .in2(_gnd_net_),
            .in3(N__37959),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_15_13_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_15_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__45315),
            .in2(_gnd_net_),
            .in3(N__37956),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_15_13_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_15_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__40257),
            .in2(_gnd_net_),
            .in3(N__37953),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_15_13_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_15_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__40232),
            .in2(_gnd_net_),
            .in3(N__37950),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_15_13_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_15_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(N__40196),
            .in2(_gnd_net_),
            .in3(N__37947),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_15_14_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_15_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__40175),
            .in2(_gnd_net_),
            .in3(N__37944),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_15_14_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_15_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__40154),
            .in2(_gnd_net_),
            .in3(N__37998),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_15_14_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_15_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__40133),
            .in2(_gnd_net_),
            .in3(N__37995),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_15_14_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_15_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__40484),
            .in2(_gnd_net_),
            .in3(N__37992),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_15_14_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_15_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__40464),
            .in2(_gnd_net_),
            .in3(N__37989),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_15_14_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_15_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__40431),
            .in2(_gnd_net_),
            .in3(N__37986),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_15_14_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_15_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__40395),
            .in2(_gnd_net_),
            .in3(N__37983),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_15_14_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_15_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__40367),
            .in2(_gnd_net_),
            .in3(N__37974),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_15_15_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_15_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__40340),
            .in2(_gnd_net_),
            .in3(N__37971),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_15_15_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_15_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__40316),
            .in2(_gnd_net_),
            .in3(N__37968),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_15_15_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_15_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__41114),
            .in2(_gnd_net_),
            .in3(N__38085),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_16_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_16_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_16_0  (
            .in0(N__45738),
            .in1(N__45416),
            .in2(N__45558),
            .in3(N__38082),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(),
            .sr(N__46863));
    defparam \delay_measurement_inst.delay_tr_reg_14_LC_15_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_14_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_14_LC_15_16_1 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_14_LC_15_16_1  (
            .in0(N__39698),
            .in1(N__38076),
            .in2(N__42902),
            .in3(N__39614),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(),
            .sr(N__46863));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_16_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_16_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_16_2  (
            .in0(N__45739),
            .in1(N__45417),
            .in2(N__45559),
            .in3(N__38040),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(),
            .sr(N__46863));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_16_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_16_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_16_3  (
            .in0(N__45414),
            .in1(N__45513),
            .in2(N__45752),
            .in3(N__38034),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(),
            .sr(N__46863));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_16_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_16_4 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_16_4  (
            .in0(N__45740),
            .in1(N__38025),
            .in2(N__45560),
            .in3(N__45419),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(),
            .sr(N__46863));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_16_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_16_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_16_5  (
            .in0(N__45415),
            .in1(N__45517),
            .in2(N__45753),
            .in3(N__38016),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(),
            .sr(N__46863));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_16_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_16_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_16_6  (
            .in0(N__45741),
            .in1(N__45418),
            .in2(N__45561),
            .in3(N__38007),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(),
            .sr(N__46863));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_17_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_17_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_17_1  (
            .in0(N__39534),
            .in1(N__39797),
            .in2(_gnd_net_),
            .in3(N__41074),
            .lcout(),
            .ltout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_17_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_17_2 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_17_2  (
            .in0(N__45443),
            .in1(N__45569),
            .in2(N__38115),
            .in3(N__45734),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47343),
            .ce(),
            .sr(N__46874));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_17_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_17_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_17_5  (
            .in0(N__45732),
            .in1(N__45444),
            .in2(N__45591),
            .in3(N__38112),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47343),
            .ce(),
            .sr(N__46874));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_17_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_17_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_17_6  (
            .in0(N__45442),
            .in1(N__45565),
            .in2(N__45751),
            .in3(N__38103),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47343),
            .ce(),
            .sr(N__46874));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_17_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_17_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_17_7  (
            .in0(N__45733),
            .in1(N__45445),
            .in2(N__45592),
            .in3(N__38094),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47343),
            .ce(),
            .sr(N__46874));
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_15_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_15_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_15_18_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_5_LC_15_18_0  (
            .in0(N__42799),
            .in1(N__43340),
            .in2(N__46336),
            .in3(N__42752),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__43380),
            .sr(N__46883));
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_15_18_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_15_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_15_18_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_8_LC_15_18_2  (
            .in0(N__42751),
            .in1(N__39575),
            .in2(_gnd_net_),
            .in3(N__43341),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__43380),
            .sr(N__46883));
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_15_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_15_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_15_18_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_3_LC_15_18_3  (
            .in0(N__40047),
            .in1(N__40010),
            .in2(_gnd_net_),
            .in3(N__46157),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__43380),
            .sr(N__46883));
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_15_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_15_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_15_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_15_LC_15_18_4  (
            .in0(N__43251),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43342),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__43380),
            .sr(N__46883));
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_15_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_15_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_15_18_5 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_14_LC_15_18_5  (
            .in0(N__43339),
            .in1(N__43252),
            .in2(_gnd_net_),
            .in3(N__42901),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__43380),
            .sr(N__46883));
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_15_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_15_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_15_18_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_1_LC_15_18_6  (
            .in0(N__46158),
            .in1(N__40083),
            .in2(N__40073),
            .in3(N__40045),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__43380),
            .sr(N__46883));
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_15_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_15_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_15_18_7 .LUT_INIT=16'b1000000010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_2_LC_15_18_7  (
            .in0(N__40046),
            .in1(N__40102),
            .in2(N__40019),
            .in3(N__46156),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__43380),
            .sr(N__46883));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_19_0  (
            .in0(N__39939),
            .in1(N__38281),
            .in2(_gnd_net_),
            .in3(N__38265),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__47329),
            .ce(N__38732),
            .sr(N__46890));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_19_1  (
            .in0(N__39935),
            .in1(N__38254),
            .in2(_gnd_net_),
            .in3(N__38238),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__47329),
            .ce(N__38732),
            .sr(N__46890));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_19_2  (
            .in0(N__39940),
            .in1(N__38233),
            .in2(_gnd_net_),
            .in3(N__38214),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__47329),
            .ce(N__38732),
            .sr(N__46890));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_19_3  (
            .in0(N__39936),
            .in1(N__38209),
            .in2(_gnd_net_),
            .in3(N__38190),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__47329),
            .ce(N__38732),
            .sr(N__46890));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_19_4  (
            .in0(N__39941),
            .in1(N__38185),
            .in2(_gnd_net_),
            .in3(N__38166),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__47329),
            .ce(N__38732),
            .sr(N__46890));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_19_5  (
            .in0(N__39937),
            .in1(N__38161),
            .in2(_gnd_net_),
            .in3(N__38142),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__47329),
            .ce(N__38732),
            .sr(N__46890));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_19_6  (
            .in0(N__39942),
            .in1(N__38137),
            .in2(_gnd_net_),
            .in3(N__38118),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__47329),
            .ce(N__38732),
            .sr(N__46890));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_19_7  (
            .in0(N__39938),
            .in1(N__38503),
            .in2(_gnd_net_),
            .in3(N__38484),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__47329),
            .ce(N__38732),
            .sr(N__46890));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_20_0  (
            .in0(N__39930),
            .in1(N__38479),
            .in2(_gnd_net_),
            .in3(N__38460),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__47325),
            .ce(N__38724),
            .sr(N__46904));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_20_1  (
            .in0(N__39889),
            .in1(N__38455),
            .in2(_gnd_net_),
            .in3(N__38436),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__47325),
            .ce(N__38724),
            .sr(N__46904));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_20_2  (
            .in0(N__39927),
            .in1(N__38431),
            .in2(_gnd_net_),
            .in3(N__38412),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__47325),
            .ce(N__38724),
            .sr(N__46904));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_20_3  (
            .in0(N__39886),
            .in1(N__38407),
            .in2(_gnd_net_),
            .in3(N__38388),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__47325),
            .ce(N__38724),
            .sr(N__46904));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_20_4  (
            .in0(N__39928),
            .in1(N__38383),
            .in2(_gnd_net_),
            .in3(N__38364),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__47325),
            .ce(N__38724),
            .sr(N__46904));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_20_5  (
            .in0(N__39887),
            .in1(N__38359),
            .in2(_gnd_net_),
            .in3(N__38340),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__47325),
            .ce(N__38724),
            .sr(N__46904));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_20_6  (
            .in0(N__39929),
            .in1(N__38335),
            .in2(_gnd_net_),
            .in3(N__38316),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__47325),
            .ce(N__38724),
            .sr(N__46904));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_20_7  (
            .in0(N__39888),
            .in1(N__38311),
            .in2(_gnd_net_),
            .in3(N__38292),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__47325),
            .ce(N__38724),
            .sr(N__46904));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_21_0  (
            .in0(N__39931),
            .in1(N__38695),
            .in2(_gnd_net_),
            .in3(N__38676),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__47321),
            .ce(N__38739),
            .sr(N__46911));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_21_1  (
            .in0(N__39923),
            .in1(N__38671),
            .in2(_gnd_net_),
            .in3(N__38652),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__47321),
            .ce(N__38739),
            .sr(N__46911));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_21_2  (
            .in0(N__39932),
            .in1(N__38647),
            .in2(_gnd_net_),
            .in3(N__38628),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__47321),
            .ce(N__38739),
            .sr(N__46911));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_21_3  (
            .in0(N__39924),
            .in1(N__38623),
            .in2(_gnd_net_),
            .in3(N__38604),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__47321),
            .ce(N__38739),
            .sr(N__46911));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_21_4  (
            .in0(N__39933),
            .in1(N__38599),
            .in2(_gnd_net_),
            .in3(N__38580),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__47321),
            .ce(N__38739),
            .sr(N__46911));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_21_5  (
            .in0(N__39925),
            .in1(N__38575),
            .in2(_gnd_net_),
            .in3(N__38556),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__47321),
            .ce(N__38739),
            .sr(N__46911));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_21_6  (
            .in0(N__39934),
            .in1(N__38551),
            .in2(_gnd_net_),
            .in3(N__38532),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__47321),
            .ce(N__38739),
            .sr(N__46911));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_21_7  (
            .in0(N__39926),
            .in1(N__38527),
            .in2(_gnd_net_),
            .in3(N__38508),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__47321),
            .ce(N__38739),
            .sr(N__46911));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_22_0  (
            .in0(N__39917),
            .in1(N__38869),
            .in2(_gnd_net_),
            .in3(N__38850),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__47318),
            .ce(N__38731),
            .sr(N__46917));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_22_1  (
            .in0(N__39921),
            .in1(N__38845),
            .in2(_gnd_net_),
            .in3(N__38826),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__47318),
            .ce(N__38731),
            .sr(N__46917));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_22_2  (
            .in0(N__39918),
            .in1(N__38821),
            .in2(_gnd_net_),
            .in3(N__38802),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__47318),
            .ce(N__38731),
            .sr(N__46917));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_22_3  (
            .in0(N__39922),
            .in1(N__38797),
            .in2(_gnd_net_),
            .in3(N__38778),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__47318),
            .ce(N__38731),
            .sr(N__46917));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_22_4  (
            .in0(N__39919),
            .in1(N__38774),
            .in2(_gnd_net_),
            .in3(N__38760),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__47318),
            .ce(N__38731),
            .sr(N__46917));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_22_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_22_5  (
            .in0(N__38753),
            .in1(N__39920),
            .in2(_gnd_net_),
            .in3(N__38757),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47318),
            .ce(N__38731),
            .sr(N__46917));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_16_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_16_6_2 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_16_6_2  (
            .in0(N__38925),
            .in1(N__38907),
            .in2(N__39099),
            .in3(N__39222),
            .lcout(\delay_measurement_inst.un1_elapsed_time_hc ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_16_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_16_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_16_7_5  (
            .in0(N__41335),
            .in1(N__41362),
            .in2(N__41285),
            .in3(N__41378),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_16_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_16_8_0 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_16_8_0  (
            .in0(N__41182),
            .in1(N__41145),
            .in2(N__41258),
            .in3(N__41212),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_16_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_16_8_1 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_16_8_1  (
            .in0(N__41705),
            .in1(N__41336),
            .in2(N__41609),
            .in3(N__41363),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH2S1_14_LC_16_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH2S1_14_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH2S1_14_LC_16_8_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH2S1_14_LC_16_8_2  (
            .in0(N__41464),
            .in1(_gnd_net_),
            .in2(N__38937),
            .in3(N__41491),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_16_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_16_8_3 .LUT_INIT=16'b0000000001011101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_16_8_3  (
            .in0(N__41492),
            .in1(N__39078),
            .in2(N__38934),
            .in3(N__41465),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_16_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_16_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_16_8_4  (
            .in0(N__41181),
            .in1(N__41579),
            .in2(N__41549),
            .in3(N__41213),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_16_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_16_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_16_8_5  (
            .in0(N__38898),
            .in1(N__39066),
            .in2(N__38916),
            .in3(N__38913),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_16_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_16_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_16_8_6  (
            .in0(N__41250),
            .in1(N__41518),
            .in2(N__41150),
            .in3(N__41429),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_16_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_16_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_16_8_7  (
            .in0(N__41211),
            .in1(N__41180),
            .in2(N__41257),
            .in3(N__41463),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_16_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_16_9_0 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_16_9_0  (
            .in0(N__39060),
            .in1(N__41462),
            .in2(N__41149),
            .in3(N__38892),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_16_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_16_9_1 .LUT_INIT=16'b0111001100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_16_9_1  (
            .in0(N__38883),
            .in1(N__39077),
            .in2(N__38874),
            .in3(N__39084),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_9_2  (
            .in0(N__41725),
            .in1(N__41404),
            .in2(N__41704),
            .in3(N__41428),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_16_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_16_9_3 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_16_9_3  (
            .in0(N__41461),
            .in1(_gnd_net_),
            .in2(N__39087),
            .in3(N__41490),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_9_4  (
            .in0(N__41542),
            .in1(N__41572),
            .in2(N__41522),
            .in3(N__41602),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_16_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_16_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_16_9_5  (
            .in0(N__41405),
            .in1(N__41281),
            .in2(N__41312),
            .in3(N__41726),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_9_6  (
            .in0(N__41210),
            .in1(N__41305),
            .in2(N__41186),
            .in3(N__41460),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI339G_25_LC_16_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI339G_25_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI339G_25_LC_16_10_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI339G_25_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__41957),
            .in2(_gnd_net_),
            .in3(N__41630),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_27_LC_16_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_27_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_27_LC_16_10_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_27_LC_16_10_1  (
            .in0(N__41934),
            .in1(N__41943),
            .in2(N__39054),
            .in3(N__38943),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7L2RA_20_LC_16_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7L2RA_20_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7L2RA_20_LC_16_10_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7L2RA_20_LC_16_10_2  (
            .in0(N__41675),
            .in1(N__39051),
            .in2(N__39045),
            .in3(N__46097),
            .lcout(\delay_measurement_inst.delay_hc_reg3lt31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_10_5  (
            .in0(N__41925),
            .in1(N__41646),
            .in2(N__41916),
            .in3(N__41655),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_16_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_16_10_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_16_10_7  (
            .in0(N__46098),
            .in1(N__41676),
            .in2(N__41798),
            .in3(N__39228),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_11_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39213),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_11_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__39192),
            .in2(N__39204),
            .in3(N__44152),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_11_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_11_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_11_2  (
            .in0(N__44135),
            .in1(N__39174),
            .in2(N__39186),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_11_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__39156),
            .in2(N__39168),
            .in3(N__44099),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_11_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__39141),
            .in2(N__39150),
            .in3(N__44063),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_11_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_11_5  (
            .in0(N__44042),
            .in1(N__39123),
            .in2(N__39135),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_11_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__39105),
            .in2(N__39117),
            .in3(N__44018),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_11_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_11_7  (
            .in0(N__44573),
            .in1(N__39363),
            .in2(N__39372),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_12_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__39348),
            .in2(N__39357),
            .in3(N__44546),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_12_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__39330),
            .in2(N__39342),
            .in3(N__44525),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_12_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_12_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_12_2  (
            .in0(N__44504),
            .in1(N__39312),
            .in2(N__39324),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_12_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__39288),
            .in2(N__39306),
            .in3(N__44480),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_12_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(N__39267),
            .in2(N__39282),
            .in3(N__44453),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_12_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__39261),
            .in2(N__39255),
            .in3(N__44423),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_12_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(N__39234),
            .in2(N__39246),
            .in3(N__44390),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_12_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(N__39471),
            .in2(N__39480),
            .in3(N__45005),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_13_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__39453),
            .in2(N__39465),
            .in3(N__44981),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_13_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__39432),
            .in2(N__39447),
            .in3(N__44960),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_13_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__39411),
            .in2(N__39426),
            .in3(N__44936),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_13_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__39390),
            .in2(N__39405),
            .in3(N__44915),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39384),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_13_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_13_5 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__44647),
            .in2(N__39381),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_13_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_13_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_13_6  (
            .in0(N__44648),
            .in1(N__44607),
            .in2(_gnd_net_),
            .in3(N__44156),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_16_14_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_16_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_16_14_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_7_LC_16_14_0  (
            .in0(N__45406),
            .in1(N__45574),
            .in2(N__45748),
            .in3(N__39558),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47375),
            .ce(),
            .sr(N__46843));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_16_14_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_16_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_16_14_1 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_8_LC_16_14_1  (
            .in0(N__45575),
            .in1(N__45716),
            .in2(N__45441),
            .in3(N__39552),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47375),
            .ce(),
            .sr(N__46843));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_16_14_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_16_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_16_14_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_9_LC_16_14_2  (
            .in0(N__45407),
            .in1(N__45576),
            .in2(N__45749),
            .in3(N__39546),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47375),
            .ce(),
            .sr(N__46843));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_14_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__39529),
            .in2(_gnd_net_),
            .in3(N__41072),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_16_14_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_16_14_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_16_14_5  (
            .in0(N__45573),
            .in1(N__45715),
            .in2(_gnd_net_),
            .in3(N__45405),
            .lcout(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_16_14_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_16_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__39530),
            .in2(_gnd_net_),
            .in3(N__41073),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_16_15_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_16_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_16_15_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_12_LC_16_15_0  (
            .in0(N__45446),
            .in1(N__45583),
            .in2(N__45750),
            .in3(N__39498),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47367),
            .ce(),
            .sr(N__46846));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_16_15_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_16_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_16_15_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_18_LC_16_15_1  (
            .in0(N__45726),
            .in1(N__45449),
            .in2(N__45598),
            .in3(N__39492),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47367),
            .ce(),
            .sr(N__46846));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_16_15_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_16_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_16_15_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_10_LC_16_15_3  (
            .in0(N__45724),
            .in1(N__45447),
            .in2(N__45596),
            .in3(N__39486),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47367),
            .ce(),
            .sr(N__46846));
    defparam \delay_measurement_inst.delay_tr_reg_15_LC_16_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_15_LC_16_15_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_15_LC_16_15_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_15_LC_16_15_4  (
            .in0(N__39699),
            .in1(N__39675),
            .in2(N__43253),
            .in3(N__39618),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47367),
            .ce(),
            .sr(N__46846));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_16_15_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_16_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_16_15_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_11_LC_16_15_5  (
            .in0(N__45725),
            .in1(N__45448),
            .in2(N__45597),
            .in3(N__39591),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47367),
            .ce(),
            .sr(N__46846));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_15_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_15_7  (
            .in0(N__47742),
            .in1(N__47605),
            .in2(N__47899),
            .in3(N__45108),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47367),
            .ce(),
            .sr(N__46846));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_16_0 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_16_16_0  (
            .in0(N__40113),
            .in1(N__46155),
            .in2(N__40020),
            .in3(N__40053),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47359),
            .ce(N__43067),
            .sr(N__46854));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_16_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_16_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_16_16_1 .LUT_INIT=16'b0100010001000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_16_16_1  (
            .in0(N__42823),
            .in1(N__42857),
            .in2(N__42783),
            .in3(N__43331),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47359),
            .ce(N__43067),
            .sr(N__46854));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_16_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_16_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_16_16_2 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_16_16_2  (
            .in0(N__42781),
            .in1(N__46308),
            .in2(N__43343),
            .in3(N__42821),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47359),
            .ce(N__43067),
            .sr(N__46854));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_16_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_16_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_16_16_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_16_16_3  (
            .in0(N__42777),
            .in1(N__42507),
            .in2(_gnd_net_),
            .in3(N__43332),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47359),
            .ce(N__43067),
            .sr(N__46854));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_16_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_16_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_16_16_4 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__42776),
            .in2(N__43344),
            .in3(N__39585),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47359),
            .ce(N__43067),
            .sr(N__46854));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_16_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_16_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_16_16_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_16_16_5  (
            .in0(N__42822),
            .in1(N__43330),
            .in2(N__46344),
            .in3(N__42782),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47359),
            .ce(N__43067),
            .sr(N__46854));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_16_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_16_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_16_16_6 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_16_16_6  (
            .in0(N__43329),
            .in1(N__42894),
            .in2(_gnd_net_),
            .in3(N__43235),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47359),
            .ce(N__43067),
            .sr(N__46854));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_16_7 .LUT_INIT=16'b1111001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_16_16_7  (
            .in0(N__43234),
            .in1(N__43148),
            .in2(N__46260),
            .in3(N__46194),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47359),
            .ce(N__43067),
            .sr(N__46854));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_16_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_16_17_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__40014),
            .in2(_gnd_net_),
            .in3(N__40112),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_17_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_16_17_2  (
            .in0(N__46147),
            .in1(N__40077),
            .in2(N__40056),
            .in3(N__40048),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47353),
            .ce(N__43062),
            .sr(N__46864));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_16_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_16_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_16_17_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_16_17_3  (
            .in0(N__40049),
            .in1(N__40015),
            .in2(_gnd_net_),
            .in3(N__46146),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47353),
            .ce(N__43062),
            .sr(N__46864));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39977),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__39777),
            .in2(N__39810),
            .in3(N__39793),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__39744),
            .in2(N__39771),
            .in3(N__39761),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_18_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_18_2  (
            .in0(N__39734),
            .in1(N__39705),
            .in2(N__39717),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_18_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_18_3  (
            .in0(N__40295),
            .in1(N__40278),
            .in2(N__42519),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__40263),
            .in2(N__40272),
            .in3(N__45314),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_18_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_18_5  (
            .in0(N__40253),
            .in1(N__40239),
            .in2(N__42711),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_18_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_18_6  (
            .in0(N__40233),
            .in1(N__40218),
            .in2(N__42477),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__40182),
            .in2(N__40212),
            .in3(N__40200),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__40161),
            .in2(N__43398),
            .in3(N__40176),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__40140),
            .in2(N__42693),
            .in3(N__40155),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__40119),
            .in2(N__42657),
            .in3(N__40134),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_19_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__40470),
            .in2(N__42624),
            .in3(N__40485),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_19_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__40446),
            .in2(N__42579),
            .in3(N__40463),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_19_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__40413),
            .in2(N__40440),
            .in3(N__40427),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_19_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__40377),
            .in2(N__40407),
            .in3(N__40391),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_19_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_19_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_19_7  (
            .in0(N__40371),
            .in1(N__42864),
            .in2(N__40353),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_20_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__40326),
            .in2(N__41040),
            .in3(N__40344),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_20_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(N__40302),
            .in2(N__41031),
            .in3(N__40320),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_20_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__41100),
            .in2(N__41022),
            .in3(N__41118),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41094),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_16_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_16_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_16_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_17_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46472),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47330),
            .ce(N__43386),
            .sr(N__46891));
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_16_20_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_16_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_16_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_18_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46510),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47330),
            .ce(N__43386),
            .sr(N__46891));
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_16_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_16_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_16_20_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_19_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__46422),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47330),
            .ce(N__43386),
            .sr(N__46891));
    defparam SB_DFF_inst_DELAY_HC1_LC_17_3_2.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_17_3_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_17_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_17_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41013),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47457),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_17_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_17_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_17_5_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_17_5_5  (
            .in0(N__40988),
            .in1(N__40959),
            .in2(_gnd_net_),
            .in3(N__43005),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_336_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_17_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_17_6_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_17_6_0 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_2_LC_17_6_0  (
            .in0(N__40877),
            .in1(N__40741),
            .in2(N__41367),
            .in3(N__40920),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47444),
            .ce(),
            .sr(N__46802));
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_17_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_17_6_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_17_6_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_15_LC_17_6_3  (
            .in0(N__40740),
            .in1(N__41469),
            .in2(N__40540),
            .in3(N__40644),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47444),
            .ce(),
            .sr(N__46802));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42969),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47437),
            .ce(N__41747),
            .sr(N__46805));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_17_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_17_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_17_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_17_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42948),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47437),
            .ce(N__41747),
            .sr(N__46805));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__42968),
            .in2(N__42927),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47429),
            .ce(N__41748),
            .sr(N__46808));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(N__42947),
            .in2(N__43614),
            .in3(N__41292),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47429),
            .ce(N__41748),
            .sr(N__46808));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(N__42926),
            .in2(N__43590),
            .in3(N__41262),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47429),
            .ce(N__41748),
            .sr(N__46808));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__43613),
            .in2(N__43566),
            .in3(N__41223),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47429),
            .ce(N__41748),
            .sr(N__46808));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(N__43589),
            .in2(N__43542),
            .in3(N__41190),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47429),
            .ce(N__41748),
            .sr(N__46808));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(N__43565),
            .in2(N__43518),
            .in3(N__41157),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47429),
            .ce(N__41748),
            .sr(N__46808));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__43541),
            .in2(N__43494),
            .in3(N__41616),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47429),
            .ce(N__41748),
            .sr(N__46808));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(N__43517),
            .in2(N__43470),
            .in3(N__41586),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47429),
            .ce(N__41748),
            .sr(N__46808));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__43493),
            .in2(N__43446),
            .in3(N__41556),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47422),
            .ce(N__41749),
            .sr(N__46811));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__43469),
            .in2(N__43422),
            .in3(N__41526),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47422),
            .ce(N__41749),
            .sr(N__46811));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__43445),
            .in2(N__43806),
            .in3(N__41499),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47422),
            .ce(N__41749),
            .sr(N__46811));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__43421),
            .in2(N__43782),
            .in3(N__41472),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47422),
            .ce(N__41749),
            .sr(N__46811));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__43805),
            .in2(N__43758),
            .in3(N__41436),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47422),
            .ce(N__41749),
            .sr(N__46811));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(N__43781),
            .in2(N__43734),
            .in3(N__41412),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47422),
            .ce(N__41749),
            .sr(N__46811));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(N__43757),
            .in2(N__43710),
            .in3(N__41391),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47422),
            .ce(N__41749),
            .sr(N__46811));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7  (
            .in0(_gnd_net_),
            .in1(N__43733),
            .in2(N__43686),
            .in3(N__41712),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47422),
            .ce(N__41749),
            .sr(N__46811));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__43709),
            .in2(N__43662),
            .in3(N__41679),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47415),
            .ce(N__41750),
            .sr(N__46815));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__43685),
            .in2(N__43638),
            .in3(N__41664),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47415),
            .ce(N__41750),
            .sr(N__46815));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__43661),
            .in2(N__43998),
            .in3(N__41661),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47415),
            .ce(N__41750),
            .sr(N__46815));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__43637),
            .in2(N__43974),
            .in3(N__41658),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47415),
            .ce(N__41750),
            .sr(N__46815));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__43997),
            .in2(N__43950),
            .in3(N__41649),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47415),
            .ce(N__41750),
            .sr(N__46815));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__43973),
            .in2(N__43926),
            .in3(N__41640),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47415),
            .ce(N__41750),
            .sr(N__46815));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(N__43949),
            .in2(N__43902),
            .in3(N__41619),
            .lcout(\delay_measurement_inst.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47415),
            .ce(N__41750),
            .sr(N__46815));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__43925),
            .in2(N__43878),
            .in3(N__41946),
            .lcout(\delay_measurement_inst.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47415),
            .ce(N__41750),
            .sr(N__46815));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__43901),
            .in2(N__43854),
            .in3(N__41937),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47407),
            .ce(N__41751),
            .sr(N__46820));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__43877),
            .in2(N__43830),
            .in3(N__41928),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47407),
            .ce(N__41751),
            .sr(N__46820));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__43853),
            .in2(N__44367),
            .in3(N__41919),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47407),
            .ce(N__41751),
            .sr(N__46820));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__43829),
            .in2(N__44226),
            .in3(N__41907),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47407),
            .ce(N__41751),
            .sr(N__46820));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41904),
            .lcout(\delay_measurement_inst.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47407),
            .ce(N__41751),
            .sr(N__46820));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_12_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_12_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_12_0  (
            .in0(N__44752),
            .in1(N__44887),
            .in2(N__42222),
            .in3(N__44052),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47398),
            .ce(),
            .sr(N__46825));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_12_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_12_1 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_12_1  (
            .in0(N__44885),
            .in1(N__42207),
            .in2(N__44031),
            .in3(N__44758),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47398),
            .ce(),
            .sr(N__46825));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_12_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_12_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_12_2  (
            .in0(N__44753),
            .in1(N__44888),
            .in2(N__42223),
            .in3(N__44007),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47398),
            .ce(),
            .sr(N__46825));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_17_12_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_17_12_3 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_7_LC_17_12_3  (
            .in0(N__44886),
            .in1(N__42208),
            .in2(N__44562),
            .in3(N__44759),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47398),
            .ce(),
            .sr(N__46825));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_12_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_12_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_12_4  (
            .in0(N__44754),
            .in1(N__44889),
            .in2(N__42224),
            .in3(N__44535),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47398),
            .ce(),
            .sr(N__46825));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_12_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_12_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_12_5  (
            .in0(N__44883),
            .in1(N__42205),
            .in2(N__44442),
            .in3(N__44756),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47398),
            .ce(),
            .sr(N__46825));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_12_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_12_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_12_6  (
            .in0(N__44755),
            .in1(N__44890),
            .in2(N__42225),
            .in3(N__44514),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47398),
            .ce(),
            .sr(N__46825));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_12_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_12_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_12_7  (
            .in0(N__44884),
            .in1(N__42206),
            .in2(N__44994),
            .in3(N__44757),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47398),
            .ce(),
            .sr(N__46825));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_13_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_13_0 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_13_0  (
            .in0(N__44875),
            .in1(N__44493),
            .in2(N__42218),
            .in3(N__44771),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__46830));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_13_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_13_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_13_1  (
            .in0(N__44764),
            .in1(N__42176),
            .in2(N__44379),
            .in3(N__44879),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__46830));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_13_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_13_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_13_2  (
            .in0(N__44876),
            .in1(N__44768),
            .in2(N__42219),
            .in3(N__44970),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__46830));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_13_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_13_3 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_13_3  (
            .in0(N__44765),
            .in1(N__42177),
            .in2(N__44949),
            .in3(N__44880),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__46830));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_13_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_13_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_13_4  (
            .in0(N__44877),
            .in1(N__44769),
            .in2(N__42220),
            .in3(N__44925),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__46830));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_13_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_13_5 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_13_5  (
            .in0(N__44766),
            .in1(N__42178),
            .in2(N__44901),
            .in3(N__44881),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__46830));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_13_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_13_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_13_6  (
            .in0(N__44878),
            .in1(N__44770),
            .in2(N__42221),
            .in3(N__44118),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__46830));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_13_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_13_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_13_7  (
            .in0(N__44767),
            .in1(N__42179),
            .in2(N__44082),
            .in3(N__44882),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__46830));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_14_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_14_0  (
            .in0(N__47572),
            .in1(N__47892),
            .in2(N__47743),
            .in3(N__45174),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47380),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.start_timer_tr_LC_17_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_17_14_1 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_17_14_1  (
            .in0(N__42084),
            .in1(N__42071),
            .in2(N__47931),
            .in3(N__42033),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47380),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_14_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_14_2  (
            .in0(N__47571),
            .in1(N__47729),
            .in2(_gnd_net_),
            .in3(N__47891),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_17_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_17_14_3 .LUT_INIT=16'b1100110111000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_17_14_3  (
            .in0(N__45959),
            .in1(N__41997),
            .in2(N__42012),
            .in3(N__45994),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47380),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__45987),
            .in2(_gnd_net_),
            .in3(N__45958),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_14_7 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_14_7  (
            .in0(N__47730),
            .in1(N__45144),
            .in2(N__47930),
            .in3(N__47573),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47380),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_17_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_17_15_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_17_15_0  (
            .in0(N__45923),
            .in1(N__41967),
            .in2(N__41979),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_17_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_17_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__42345),
            .in2(N__42357),
            .in3(N__45119),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_17_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_17_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__42324),
            .in2(N__42339),
            .in3(N__45278),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_17_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_17_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__42309),
            .in2(N__42318),
            .in3(N__45248),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_17_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_17_15_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_17_15_4  (
            .in0(N__45221),
            .in1(N__42291),
            .in2(N__42303),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_17_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_17_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__42276),
            .in2(N__42285),
            .in3(N__46070),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_17_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_17_15_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_17_15_6  (
            .in0(N__46043),
            .in1(N__42258),
            .in2(N__42270),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_17_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_17_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__42252),
            .in2(N__42240),
            .in3(N__45077),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_17_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_17_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__42456),
            .in2(N__42465),
            .in3(N__45044),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_17_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_17_16_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_17_16_1  (
            .in0(N__46013),
            .in1(N__42450),
            .in2(N__43083),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_17_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_17_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__42432),
            .in2(N__42444),
            .in3(N__45890),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_17_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_17_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__42414),
            .in2(N__42426),
            .in3(N__45863),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_17_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_17_16_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_17_16_4  (
            .in0(N__45833),
            .in1(N__42393),
            .in2(N__42408),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_17_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_17_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__42375),
            .in2(N__42387),
            .in3(N__47957),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_17_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_17_16_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_17_16_6  (
            .in0(N__47480),
            .in1(N__42369),
            .in2(N__43188),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_17_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_17_16_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_17_16_7  (
            .in0(N__45189),
            .in1(N__42363),
            .in2(N__43173),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_17_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_17_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__42567),
            .in2(N__42546),
            .in3(N__45161),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_17_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_17_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__42561),
            .in2(N__42537),
            .in3(N__45794),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_17_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_17_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__42555),
            .in2(N__42528),
            .in3(N__45776),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_17_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_17_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42549),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_17_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_17_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_17_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46473),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__43063),
            .sr(N__46855));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_17_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_17_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_17_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46515),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__43063),
            .sr(N__46855));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_17_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_17_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_17_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46433),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__43063),
            .sr(N__46855));
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_17_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_17_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_17_18_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_4_LC_17_18_0  (
            .in0(N__42773),
            .in1(N__43301),
            .in2(N__46307),
            .in3(N__42824),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47354),
            .ce(N__43384),
            .sr(N__46865));
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_17_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_17_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_17_18_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_7_LC_17_18_1  (
            .in0(N__43300),
            .in1(N__42506),
            .in2(_gnd_net_),
            .in3(N__42774),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47354),
            .ce(N__43384),
            .sr(N__46865));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_17_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_17_18_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__43239),
            .in2(_gnd_net_),
            .in3(N__42903),
            .lcout(\phase_controller_inst1.stoper_tr.N_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_17_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_17_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_17_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_16_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46383),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47354),
            .ce(N__43384),
            .sr(N__46865));
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_17_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_17_19_0 .LUT_INIT=16'b0000110000001101;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_6_LC_17_19_0  (
            .in0(N__43299),
            .in1(N__42858),
            .in2(N__42828),
            .in3(N__42775),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47344),
            .ce(N__43385),
            .sr(N__46875));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_17_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_17_19_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_17_19_1  (
            .in0(N__46471),
            .in1(N__46381),
            .in2(N__46432),
            .in3(N__46506),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_17_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_17_19_2 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42699),
            .in3(N__46272),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_17_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_17_19_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_10_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42696),
            .in3(N__43109),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47344),
            .ce(N__43385),
            .sr(N__46875));
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_17_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_17_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_17_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_11_LC_17_19_4  (
            .in0(N__43137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42681),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47344),
            .ce(N__43385),
            .sr(N__46875));
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_17_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_17_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_17_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_12_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__43138),
            .in2(_gnd_net_),
            .in3(N__42648),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47344),
            .ce(N__43385),
            .sr(N__46875));
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_17_19_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_17_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_17_19_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_13_LC_17_19_6  (
            .in0(N__43139),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42607),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47344),
            .ce(N__43385),
            .sr(N__46875));
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_17_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_17_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_17_19_7 .LUT_INIT=16'b1011101010111011;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_9_LC_17_19_7  (
            .in0(N__46256),
            .in1(N__43140),
            .in2(N__43260),
            .in3(N__46193),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47344),
            .ce(N__43385),
            .sr(N__46875));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_20_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__43302),
            .in2(_gnd_net_),
            .in3(N__43257),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47336),
            .ce(N__43068),
            .sr(N__46884));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_17_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_17_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_17_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46382),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47336),
            .ce(N__43068),
            .sr(N__46884));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_17_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_17_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_17_20_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(N__43141),
            .in2(_gnd_net_),
            .in3(N__43110),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47336),
            .ce(N__43068),
            .sr(N__46884));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43001),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0  (
            .in0(N__44320),
            .in1(N__42967),
            .in2(_gnd_net_),
            .in3(N__42951),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__47445),
            .ce(N__44205),
            .sr(N__46803));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1  (
            .in0(N__44342),
            .in1(N__42946),
            .in2(_gnd_net_),
            .in3(N__42930),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__47445),
            .ce(N__44205),
            .sr(N__46803));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2  (
            .in0(N__44321),
            .in1(N__42925),
            .in2(_gnd_net_),
            .in3(N__42906),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__47445),
            .ce(N__44205),
            .sr(N__46803));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3  (
            .in0(N__44343),
            .in1(N__43612),
            .in2(_gnd_net_),
            .in3(N__43593),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__47445),
            .ce(N__44205),
            .sr(N__46803));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4  (
            .in0(N__44322),
            .in1(N__43588),
            .in2(_gnd_net_),
            .in3(N__43569),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__47445),
            .ce(N__44205),
            .sr(N__46803));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5  (
            .in0(N__44344),
            .in1(N__43564),
            .in2(_gnd_net_),
            .in3(N__43545),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__47445),
            .ce(N__44205),
            .sr(N__46803));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6  (
            .in0(N__44323),
            .in1(N__43540),
            .in2(_gnd_net_),
            .in3(N__43521),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__47445),
            .ce(N__44205),
            .sr(N__46803));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7  (
            .in0(N__44345),
            .in1(N__43516),
            .in2(_gnd_net_),
            .in3(N__43497),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__47445),
            .ce(N__44205),
            .sr(N__46803));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0  (
            .in0(N__44333),
            .in1(N__43492),
            .in2(_gnd_net_),
            .in3(N__43473),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__47438),
            .ce(N__44207),
            .sr(N__46806));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1  (
            .in0(N__44349),
            .in1(N__43468),
            .in2(_gnd_net_),
            .in3(N__43449),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__47438),
            .ce(N__44207),
            .sr(N__46806));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2  (
            .in0(N__44330),
            .in1(N__43444),
            .in2(_gnd_net_),
            .in3(N__43425),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__47438),
            .ce(N__44207),
            .sr(N__46806));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3  (
            .in0(N__44346),
            .in1(N__43420),
            .in2(_gnd_net_),
            .in3(N__43401),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__47438),
            .ce(N__44207),
            .sr(N__46806));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4  (
            .in0(N__44331),
            .in1(N__43804),
            .in2(_gnd_net_),
            .in3(N__43785),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__47438),
            .ce(N__44207),
            .sr(N__46806));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5  (
            .in0(N__44347),
            .in1(N__43780),
            .in2(_gnd_net_),
            .in3(N__43761),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__47438),
            .ce(N__44207),
            .sr(N__46806));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6  (
            .in0(N__44332),
            .in1(N__43756),
            .in2(_gnd_net_),
            .in3(N__43737),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__47438),
            .ce(N__44207),
            .sr(N__46806));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7  (
            .in0(N__44348),
            .in1(N__43732),
            .in2(_gnd_net_),
            .in3(N__43713),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__47438),
            .ce(N__44207),
            .sr(N__46806));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0  (
            .in0(N__44334),
            .in1(N__43708),
            .in2(_gnd_net_),
            .in3(N__43689),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_18_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__47430),
            .ce(N__44206),
            .sr(N__46809));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1  (
            .in0(N__44338),
            .in1(N__43684),
            .in2(_gnd_net_),
            .in3(N__43665),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__47430),
            .ce(N__44206),
            .sr(N__46809));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2  (
            .in0(N__44335),
            .in1(N__43660),
            .in2(_gnd_net_),
            .in3(N__43641),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__47430),
            .ce(N__44206),
            .sr(N__46809));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3  (
            .in0(N__44339),
            .in1(N__43636),
            .in2(_gnd_net_),
            .in3(N__43617),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__47430),
            .ce(N__44206),
            .sr(N__46809));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4  (
            .in0(N__44336),
            .in1(N__43996),
            .in2(_gnd_net_),
            .in3(N__43977),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__47430),
            .ce(N__44206),
            .sr(N__46809));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5  (
            .in0(N__44340),
            .in1(N__43972),
            .in2(_gnd_net_),
            .in3(N__43953),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__47430),
            .ce(N__44206),
            .sr(N__46809));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6  (
            .in0(N__44337),
            .in1(N__43948),
            .in2(_gnd_net_),
            .in3(N__43929),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__47430),
            .ce(N__44206),
            .sr(N__46809));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7  (
            .in0(N__44341),
            .in1(N__43924),
            .in2(_gnd_net_),
            .in3(N__43905),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__47430),
            .ce(N__44206),
            .sr(N__46809));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0  (
            .in0(N__44324),
            .in1(N__43900),
            .in2(_gnd_net_),
            .in3(N__43881),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__47423),
            .ce(N__44211),
            .sr(N__46812));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1  (
            .in0(N__44328),
            .in1(N__43876),
            .in2(_gnd_net_),
            .in3(N__43857),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__47423),
            .ce(N__44211),
            .sr(N__46812));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2  (
            .in0(N__44325),
            .in1(N__43852),
            .in2(_gnd_net_),
            .in3(N__43833),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__47423),
            .ce(N__44211),
            .sr(N__46812));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3  (
            .in0(N__44329),
            .in1(N__43828),
            .in2(_gnd_net_),
            .in3(N__43809),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__47423),
            .ce(N__44211),
            .sr(N__46812));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4  (
            .in0(N__44326),
            .in1(N__44366),
            .in2(_gnd_net_),
            .in3(N__44352),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__47423),
            .ce(N__44211),
            .sr(N__46812));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5  (
            .in0(N__44225),
            .in1(N__44327),
            .in2(_gnd_net_),
            .in3(N__44229),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47423),
            .ce(N__44211),
            .sr(N__46812));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_11_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__44175),
            .in2(N__44163),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_11_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_11_1  (
            .in0(_gnd_net_),
            .in1(N__44136),
            .in2(_gnd_net_),
            .in3(N__44106),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_11_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__44583),
            .in2(N__44103),
            .in3(N__44067),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_11_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(N__44064),
            .in2(_gnd_net_),
            .in3(N__44046),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_11_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__44043),
            .in2(_gnd_net_),
            .in3(N__44022),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_11_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__44019),
            .in2(_gnd_net_),
            .in3(N__44001),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_11_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__44574),
            .in2(_gnd_net_),
            .in3(N__44550),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_11_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(N__44547),
            .in2(_gnd_net_),
            .in3(N__44529),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_12_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__44526),
            .in2(_gnd_net_),
            .in3(N__44508),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_12_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__44505),
            .in2(_gnd_net_),
            .in3(N__44487),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_12_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_12_2  (
            .in0(_gnd_net_),
            .in1(N__44484),
            .in2(_gnd_net_),
            .in3(N__44457),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_12_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_12_3  (
            .in0(_gnd_net_),
            .in1(N__44454),
            .in2(_gnd_net_),
            .in3(N__44430),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_12_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_12_4  (
            .in0(_gnd_net_),
            .in1(N__44427),
            .in2(_gnd_net_),
            .in3(N__44394),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_12_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(N__44391),
            .in2(_gnd_net_),
            .in3(N__44370),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_12_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(N__45006),
            .in2(_gnd_net_),
            .in3(N__44985),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_12_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_12_7  (
            .in0(_gnd_net_),
            .in1(N__44982),
            .in2(_gnd_net_),
            .in3(N__44964),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_13_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__44961),
            .in2(_gnd_net_),
            .in3(N__44940),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_13_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__44937),
            .in2(_gnd_net_),
            .in3(N__44919),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_13_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_13_2  (
            .in0(_gnd_net_),
            .in1(N__44916),
            .in2(_gnd_net_),
            .in3(N__44904),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_18_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_18_13_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__47734),
            .in2(_gnd_net_),
            .in3(N__47536),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_18_13_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_18_13_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__44874),
            .in2(_gnd_net_),
            .in3(N__44763),
            .lcout(\phase_controller_slave.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_18_13_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_18_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(N__44643),
            .in2(_gnd_net_),
            .in3(N__44611),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__45132),
            .in2(N__45927),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__45126),
            .in2(_gnd_net_),
            .in3(N__45096),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__45813),
            .in2(N__45282),
            .in3(N__45093),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__45249),
            .in2(_gnd_net_),
            .in3(N__45090),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__45222),
            .in2(_gnd_net_),
            .in3(N__45087),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__46074),
            .in2(_gnd_net_),
            .in3(N__45084),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__46044),
            .in2(_gnd_net_),
            .in3(N__45081),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__45078),
            .in2(_gnd_net_),
            .in3(N__45048),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__45045),
            .in2(_gnd_net_),
            .in3(N__45009),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__46014),
            .in2(_gnd_net_),
            .in3(N__45207),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__45891),
            .in2(_gnd_net_),
            .in3(N__45204),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__45864),
            .in2(_gnd_net_),
            .in3(N__45201),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__45834),
            .in2(_gnd_net_),
            .in3(N__45198),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__47958),
            .in2(_gnd_net_),
            .in3(N__45195),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__47481),
            .in2(_gnd_net_),
            .in3(N__45192),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__45188),
            .in2(_gnd_net_),
            .in3(N__45168),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__45165),
            .in2(_gnd_net_),
            .in3(N__45135),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__45795),
            .in2(_gnd_net_),
            .in3(N__45819),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_16_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__45777),
            .in2(_gnd_net_),
            .in3(N__45816),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_18_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_18_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__45995),
            .in2(_gnd_net_),
            .in3(N__45956),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_17_0 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_17_0  (
            .in0(N__47621),
            .in1(N__47789),
            .in2(N__45804),
            .in3(N__47921),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47368),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_17_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_17_1  (
            .in0(N__47781),
            .in1(N__47624),
            .in2(N__47936),
            .in3(N__45783),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47368),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_18_17_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_18_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_18_17_2 .LUT_INIT=16'b1010101010000010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_5_LC_18_17_2  (
            .in0(N__45765),
            .in1(N__45731),
            .in2(N__45600),
            .in3(N__45450),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47368),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_17_3 .LUT_INIT=16'b1010100010001010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_17_3  (
            .in0(N__45291),
            .in1(N__47627),
            .in2(N__47790),
            .in3(N__47924),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47368),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_17_4 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_17_4  (
            .in0(N__47622),
            .in1(N__47922),
            .in2(N__45261),
            .in3(N__47784),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47368),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_17_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_17_5  (
            .in0(N__47782),
            .in1(N__47625),
            .in2(N__47937),
            .in3(N__45231),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47368),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_17_6 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_17_6  (
            .in0(N__47623),
            .in1(N__47923),
            .in2(N__46086),
            .in3(N__47785),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47368),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_17_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_17_7  (
            .in0(N__47783),
            .in1(N__47626),
            .in2(N__47938),
            .in3(N__46056),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47368),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_18_0 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_18_0  (
            .in0(N__47774),
            .in1(N__47909),
            .in2(N__47628),
            .in3(N__46026),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47361),
            .ce(),
            .sr(N__46856));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_18_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_18_18_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_18_18_1  (
            .in0(N__45999),
            .in1(N__45922),
            .in2(_gnd_net_),
            .in3(N__45957),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_18_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_18_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_18_18_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_18_18_2  (
            .in0(N__47777),
            .in1(N__47908),
            .in2(N__45930),
            .in3(N__47620),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47361),
            .ce(),
            .sr(N__46856));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_18_3 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_18_3  (
            .in0(N__45900),
            .in1(N__47778),
            .in2(N__47631),
            .in3(N__47925),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47361),
            .ce(),
            .sr(N__46856));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_18_4 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_18_4  (
            .in0(N__47775),
            .in1(N__47910),
            .in2(N__47629),
            .in3(N__45873),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47361),
            .ce(),
            .sr(N__46856));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_18_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_18_5  (
            .in0(N__47906),
            .in1(N__47779),
            .in2(N__45846),
            .in3(N__47615),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47361),
            .ce(),
            .sr(N__46856));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_18_6 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_18_6  (
            .in0(N__47776),
            .in1(N__47911),
            .in2(N__47630),
            .in3(N__47967),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47361),
            .ce(),
            .sr(N__46856));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_18_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_18_7  (
            .in0(N__47907),
            .in1(N__47780),
            .in2(N__47646),
            .in3(N__47616),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47361),
            .ce(),
            .sr(N__46856));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_18_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_18_19_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_18_19_4  (
            .in0(N__46514),
            .in1(N__46470),
            .in2(N__46434),
            .in3(N__46380),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_18_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_18_19_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_18_19_5  (
            .in0(N__46340),
            .in1(N__46306),
            .in2(N__46275),
            .in3(N__46271),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_18_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_18_19_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_18_19_6  (
            .in0(N__46248),
            .in1(N__46215),
            .in2(N__46197),
            .in3(N__46192),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_20_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_20_10_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(N__46116),
            .in2(_gnd_net_),
            .in3(N__46107),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MAIN
